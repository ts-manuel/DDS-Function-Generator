// NiosII_Processor_LCD.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module NiosII_Processor_LCD (
		input  wire        BackLight_PWM_clk_clk,                    //                 BackLight_PWM_clk.clk
		output wire [7:0]  BackLight_PWM_external_connection_export, // BackLight_PWM_external_connection.export
		input  wire        BackLight_PWM_reset_reset_n,              //               BackLight_PWM_reset.reset_n
		input  wire [1:0]  BackLight_PWM_s1_address,                 //                  BackLight_PWM_s1.address
		input  wire        BackLight_PWM_s1_write_n,                 //                                  .write_n
		input  wire [31:0] BackLight_PWM_s1_writedata,               //                                  .writedata
		input  wire        BackLight_PWM_s1_chipselect,              //                                  .chipselect
		output wire [31:0] BackLight_PWM_s1_readdata,                //                                  .readdata
		input  wire        Control_clk_clk,                          //                       Control_clk.clk
		output wire [4:0]  Control_external_connection_export,       //       Control_external_connection.export
		input  wire        Control_reset_reset_n,                    //                     Control_reset.reset_n
		input  wire [2:0]  Control_s1_address,                       //                        Control_s1.address
		input  wire        Control_s1_write_n,                       //                                  .write_n
		input  wire [31:0] Control_s1_writedata,                     //                                  .writedata
		input  wire        Control_s1_chipselect,                    //                                  .chipselect
		output wire [31:0] Control_s1_readdata,                      //                                  .readdata
		input  wire        Data_clk_clk,                             //                          Data_clk.clk
		input  wire        Data_reset_reset_n,                       //                        Data_reset.reset_n
		input  wire [1:0]  Data_s1_address,                          //                           Data_s1.address
		input  wire        Data_s1_write_n,                          //                                  .write_n
		input  wire [31:0] Data_s1_writedata,                        //                                  .writedata
		input  wire        Data_s1_chipselect,                       //                                  .chipselect
		output wire [31:0] Data_s1_readdata,                         //                                  .readdata
		output wire [7:0]  data_external_connection_export           //          data_external_connection.export
	);

	NiosII_Processor_LCD_BackLight_PWM backlight_pwm (
		.clk        (BackLight_PWM_clk_clk),                    //                 clk.clk
		.reset_n    (BackLight_PWM_reset_reset_n),              //               reset.reset_n
		.address    (BackLight_PWM_s1_address),                 //                  s1.address
		.write_n    (BackLight_PWM_s1_write_n),                 //                    .write_n
		.writedata  (BackLight_PWM_s1_writedata),               //                    .writedata
		.chipselect (BackLight_PWM_s1_chipselect),              //                    .chipselect
		.readdata   (BackLight_PWM_s1_readdata),                //                    .readdata
		.out_port   (BackLight_PWM_external_connection_export)  // external_connection.export
	);

	NiosII_Processor_LCD_Control control (
		.clk        (Control_clk_clk),                    //                 clk.clk
		.reset_n    (Control_reset_reset_n),              //               reset.reset_n
		.address    (Control_s1_address),                 //                  s1.address
		.write_n    (Control_s1_write_n),                 //                    .write_n
		.writedata  (Control_s1_writedata),               //                    .writedata
		.chipselect (Control_s1_chipselect),              //                    .chipselect
		.readdata   (Control_s1_readdata),                //                    .readdata
		.out_port   (Control_external_connection_export)  // external_connection.export
	);

	NiosII_Processor_LCD_BackLight_PWM data (
		.clk        (Data_clk_clk),                    //                 clk.clk
		.reset_n    (Data_reset_reset_n),              //               reset.reset_n
		.address    (Data_s1_address),                 //                  s1.address
		.write_n    (Data_s1_write_n),                 //                    .write_n
		.writedata  (Data_s1_writedata),               //                    .writedata
		.chipselect (Data_s1_chipselect),              //                    .chipselect
		.readdata   (Data_s1_readdata),                //                    .readdata
		.out_port   (data_external_connection_export)  // external_connection.export
	);

endmodule
