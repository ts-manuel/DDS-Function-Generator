// NiosII_Processor.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module NiosII_Processor (
		input  wire [1:0]  btn_ch_onoff_export,              //              btn_ch_onoff.export
		input  wire [5:0]  btn_display_export,               //               btn_display.export
		input  wire [4:0]  btn_encoder_export,               //               btn_encoder.export
		input  wire        clk_clk,                          //                       clk.clk
		output wire        cpu_reset,                        //                       cpu.reset
		output wire [31:0] dds0_am_modindex_export,          //          dds0_am_modindex.export
		output wire [31:0] dds0_am_modphasestep_export,      //      dds0_am_modphasestep.export
		output wire [31:0] dds0_fm_moddeviationphase_export, // dds0_fm_moddeviationphase.export
		output wire [31:0] dds0_fm_modphasestep_export,      //      dds0_fm_modphasestep.export
		output wire        dds0_outputrelay_export,          //          dds0_outputrelay.export
		output wire [31:0] dds0_phaseoffset_export,          //          dds0_phaseoffset.export
		output wire [31:0] dds0_phasestep_export,            //            dds0_phasestep.export
		output wire [31:0] dds0_pm_modindex_export,          //          dds0_pm_modindex.export
		output wire [31:0] dds0_pm_modphasestep_export,      //      dds0_pm_modphasestep.export
		output wire [15:0] dds0_pwm_amplitude_export,        //        dds0_pwm_amplitude.export
		output wire [15:0] dds0_pwm_offset_export,           //           dds0_pwm_offset.export
		output wire [31:0] dds1_am_modindex_export,          //          dds1_am_modindex.export
		output wire [31:0] dds1_am_modphasestep_export,      //      dds1_am_modphasestep.export
		output wire [31:0] dds1_fm_moddeviationphase_export, // dds1_fm_moddeviationphase.export
		output wire [31:0] dds1_fm_modphasestep_export,      //      dds1_fm_modphasestep.export
		output wire        dds1_outputrelay_export,          //          dds1_outputrelay.export
		output wire [31:0] dds1_phaseoffset_export,          //          dds1_phaseoffset.export
		output wire [31:0] dds1_phasestep_export,            //            dds1_phasestep.export
		output wire [31:0] dds1_pm_modindex_export,          //          dds1_pm_modindex.export
		output wire [31:0] dds1_pm_modphasestep_export,      //      dds1_pm_modphasestep.export
		output wire [15:0] dds1_pwm_amplitude_export,        //        dds1_pwm_amplitude.export
		output wire [15:0] dds1_pwm_offset_export,           //           dds1_pwm_offset.export
		output wire [1:0]  dds_reset_export,                 //                 dds_reset.export
		input  wire [7:0]  keypad_input_export,              //              keypad_input.export
		output wire [7:0]  lcd_backlight_pwm_export,         //         lcd_backlight_pwm.export
		output wire [4:0]  lcd_control_export,               //               lcd_control.export
		output wire [7:0]  lcd_data_export,                  //                  lcd_data.export
		output wire [4:0]  lcd_dma_address,                  //                   lcd_dma.address
		output wire        lcd_dma_chipselect,               //                          .chipselect
		input  wire        lcd_dma_waitrequest,              //                          .waitrequest
		output wire        lcd_dma_write_n,                  //                          .write_n
		output wire [7:0]  lcd_dma_writedata,                //                          .writedata
		output wire        led_debug_export,                 //                 led_debug.export
		input  wire [5:0]  lookup_ram_isr_1_export,          //          lookup_ram_isr_1.export
		input  wire [9:0]  ram_dds0_address,                 //                  ram_dds0.address
		input  wire        ram_dds0_chipselect,              //                          .chipselect
		input  wire        ram_dds0_clken,                   //                          .clken
		input  wire        ram_dds0_write,                   //                          .write
		output wire [15:0] ram_dds0_readdata,                //                          .readdata
		input  wire [15:0] ram_dds0_writedata,               //                          .writedata
		input  wire [1:0]  ram_dds0_byteenable,              //                          .byteenable
		input  wire [9:0]  ram_dds0_am_address,              //               ram_dds0_am.address
		input  wire        ram_dds0_am_chipselect,           //                          .chipselect
		input  wire        ram_dds0_am_clken,                //                          .clken
		input  wire        ram_dds0_am_write,                //                          .write
		output wire [15:0] ram_dds0_am_readdata,             //                          .readdata
		input  wire [15:0] ram_dds0_am_writedata,            //                          .writedata
		input  wire [1:0]  ram_dds0_am_byteenable,           //                          .byteenable
		input  wire        ram_dds0_clk_clk,                 //              ram_dds0_clk.clk
		input  wire [9:0]  ram_dds0_fm_address,              //               ram_dds0_fm.address
		input  wire        ram_dds0_fm_chipselect,           //                          .chipselect
		input  wire        ram_dds0_fm_clken,                //                          .clken
		input  wire        ram_dds0_fm_write,                //                          .write
		output wire [15:0] ram_dds0_fm_readdata,             //                          .readdata
		input  wire [15:0] ram_dds0_fm_writedata,            //                          .writedata
		input  wire [1:0]  ram_dds0_fm_byteenable,           //                          .byteenable
		input  wire        ram_dds0_reset_reset_n,           //            ram_dds0_reset.reset_n
		input  wire [9:0]  ram_dds1_address,                 //                  ram_dds1.address
		input  wire        ram_dds1_chipselect,              //                          .chipselect
		input  wire        ram_dds1_clken,                   //                          .clken
		input  wire        ram_dds1_write,                   //                          .write
		output wire [15:0] ram_dds1_readdata,                //                          .readdata
		input  wire [15:0] ram_dds1_writedata,               //                          .writedata
		input  wire [1:0]  ram_dds1_byteenable,              //                          .byteenable
		input  wire [9:0]  ram_dds1_am_address,              //               ram_dds1_am.address
		input  wire        ram_dds1_am_chipselect,           //                          .chipselect
		input  wire        ram_dds1_am_clken,                //                          .clken
		input  wire        ram_dds1_am_write,                //                          .write
		output wire [15:0] ram_dds1_am_readdata,             //                          .readdata
		input  wire [15:0] ram_dds1_am_writedata,            //                          .writedata
		input  wire [1:0]  ram_dds1_am_byteenable,           //                          .byteenable
		input  wire [9:0]  ram_dds1_fm_address,              //               ram_dds1_fm.address
		input  wire        ram_dds1_fm_chipselect,           //                          .chipselect
		input  wire        ram_dds1_fm_clken,                //                          .clken
		input  wire        ram_dds1_fm_write,                //                          .write
		output wire [15:0] ram_dds1_fm_readdata,             //                          .readdata
		input  wire [15:0] ram_dds1_fm_writedata,            //                          .writedata
		input  wire [1:0]  ram_dds1_fm_byteenable,           //                          .byteenable
		input  wire        sd_spi_MISO,                      //                    sd_spi.MISO
		output wire        sd_spi_MOSI,                      //                          .MOSI
		output wire        sd_spi_SCLK,                      //                          .SCLK
		output wire        sd_spi_SS_n,                      //                          .SS_n
		output wire [4:0]  spi_dma_address,                  //                   spi_dma.address
		output wire        spi_dma_chipselect,               //                          .chipselect
		output wire        spi_dma_read_n,                   //                          .read_n
		input  wire [7:0]  spi_dma_readdata,                 //                          .readdata
		input  wire        spi_dma_readdatavalid,            //                          .readdatavalid
		input  wire        spi_dma_waitrequest               //                          .waitrequest
	);

	wire         nios_cpu_debug_reset_request_reset;                        // NIOS_CPU:debug_reset_request -> rst_controller:reset_in0
	wire  [31:0] nios_cpu_data_master_readdata;                             // mm_interconnect_0:NIOS_CPU_data_master_readdata -> NIOS_CPU:d_readdata
	wire         nios_cpu_data_master_waitrequest;                          // mm_interconnect_0:NIOS_CPU_data_master_waitrequest -> NIOS_CPU:d_waitrequest
	wire         nios_cpu_data_master_debugaccess;                          // NIOS_CPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOS_CPU_data_master_debugaccess
	wire  [19:0] nios_cpu_data_master_address;                              // NIOS_CPU:d_address -> mm_interconnect_0:NIOS_CPU_data_master_address
	wire   [3:0] nios_cpu_data_master_byteenable;                           // NIOS_CPU:d_byteenable -> mm_interconnect_0:NIOS_CPU_data_master_byteenable
	wire         nios_cpu_data_master_read;                                 // NIOS_CPU:d_read -> mm_interconnect_0:NIOS_CPU_data_master_read
	wire         nios_cpu_data_master_write;                                // NIOS_CPU:d_write -> mm_interconnect_0:NIOS_CPU_data_master_write
	wire  [31:0] nios_cpu_data_master_writedata;                            // NIOS_CPU:d_writedata -> mm_interconnect_0:NIOS_CPU_data_master_writedata
	wire         lcd_dma_read_master_chipselect;                            // LCD_DMA:read_chipselect -> mm_interconnect_0:LCD_DMA_read_master_chipselect
	wire   [7:0] lcd_dma_read_master_readdata;                              // mm_interconnect_0:LCD_DMA_read_master_readdata -> LCD_DMA:read_readdata
	wire         lcd_dma_read_master_waitrequest;                           // mm_interconnect_0:LCD_DMA_read_master_waitrequest -> LCD_DMA:read_waitrequest
	wire  [14:0] lcd_dma_read_master_address;                               // LCD_DMA:read_address -> mm_interconnect_0:LCD_DMA_read_master_address
	wire         lcd_dma_read_master_read;                                  // LCD_DMA:read_read_n -> mm_interconnect_0:LCD_DMA_read_master_read
	wire         lcd_dma_read_master_readdatavalid;                         // mm_interconnect_0:LCD_DMA_read_master_readdatavalid -> LCD_DMA:read_readdatavalid
	wire         spi_dma_write_master_chipselect;                           // SPI_DMA:write_chipselect -> mm_interconnect_0:SPI_DMA_write_master_chipselect
	wire         spi_dma_write_master_waitrequest;                          // mm_interconnect_0:SPI_DMA_write_master_waitrequest -> SPI_DMA:write_waitrequest
	wire  [14:0] spi_dma_write_master_address;                              // SPI_DMA:write_address -> mm_interconnect_0:SPI_DMA_write_master_address
	wire         spi_dma_write_master_write;                                // SPI_DMA:write_write_n -> mm_interconnect_0:SPI_DMA_write_master_write
	wire   [7:0] spi_dma_write_master_writedata;                            // SPI_DMA:write_writedata -> mm_interconnect_0:SPI_DMA_write_master_writedata
	wire  [31:0] nios_cpu_instruction_master_readdata;                      // mm_interconnect_0:NIOS_CPU_instruction_master_readdata -> NIOS_CPU:i_readdata
	wire         nios_cpu_instruction_master_waitrequest;                   // mm_interconnect_0:NIOS_CPU_instruction_master_waitrequest -> NIOS_CPU:i_waitrequest
	wire  [19:0] nios_cpu_instruction_master_address;                       // NIOS_CPU:i_address -> mm_interconnect_0:NIOS_CPU_instruction_master_address
	wire         nios_cpu_instruction_master_read;                          // NIOS_CPU:i_read -> mm_interconnect_0:NIOS_CPU_instruction_master_read
	wire         mm_interconnect_0_dds0_am_modindex_s1_chipselect;          // mm_interconnect_0:DDS0_AM_ModIndex_s1_chipselect -> DDS0:AM_ModIndex_s1_chipselect
	wire  [31:0] mm_interconnect_0_dds0_am_modindex_s1_readdata;            // DDS0:AM_ModIndex_s1_readdata -> mm_interconnect_0:DDS0_AM_ModIndex_s1_readdata
	wire   [1:0] mm_interconnect_0_dds0_am_modindex_s1_address;             // mm_interconnect_0:DDS0_AM_ModIndex_s1_address -> DDS0:AM_ModIndex_s1_address
	wire         mm_interconnect_0_dds0_am_modindex_s1_write;               // mm_interconnect_0:DDS0_AM_ModIndex_s1_write -> DDS0:AM_ModIndex_s1_write_n
	wire  [31:0] mm_interconnect_0_dds0_am_modindex_s1_writedata;           // mm_interconnect_0:DDS0_AM_ModIndex_s1_writedata -> DDS0:AM_ModIndex_s1_writedata
	wire         mm_interconnect_0_dds1_am_modindex_s1_chipselect;          // mm_interconnect_0:DDS1_AM_ModIndex_s1_chipselect -> DDS1:AM_ModIndex_s1_chipselect
	wire  [31:0] mm_interconnect_0_dds1_am_modindex_s1_readdata;            // DDS1:AM_ModIndex_s1_readdata -> mm_interconnect_0:DDS1_AM_ModIndex_s1_readdata
	wire   [1:0] mm_interconnect_0_dds1_am_modindex_s1_address;             // mm_interconnect_0:DDS1_AM_ModIndex_s1_address -> DDS1:AM_ModIndex_s1_address
	wire         mm_interconnect_0_dds1_am_modindex_s1_write;               // mm_interconnect_0:DDS1_AM_ModIndex_s1_write -> DDS1:AM_ModIndex_s1_write_n
	wire  [31:0] mm_interconnect_0_dds1_am_modindex_s1_writedata;           // mm_interconnect_0:DDS1_AM_ModIndex_s1_writedata -> DDS1:AM_ModIndex_s1_writedata
	wire         mm_interconnect_0_dds0_am_modphasestep_s1_chipselect;      // mm_interconnect_0:DDS0_AM_ModPhaseStep_s1_chipselect -> DDS0:AM_ModPhaseStep_s1_chipselect
	wire  [31:0] mm_interconnect_0_dds0_am_modphasestep_s1_readdata;        // DDS0:AM_ModPhaseStep_s1_readdata -> mm_interconnect_0:DDS0_AM_ModPhaseStep_s1_readdata
	wire   [1:0] mm_interconnect_0_dds0_am_modphasestep_s1_address;         // mm_interconnect_0:DDS0_AM_ModPhaseStep_s1_address -> DDS0:AM_ModPhaseStep_s1_address
	wire         mm_interconnect_0_dds0_am_modphasestep_s1_write;           // mm_interconnect_0:DDS0_AM_ModPhaseStep_s1_write -> DDS0:AM_ModPhaseStep_s1_write_n
	wire  [31:0] mm_interconnect_0_dds0_am_modphasestep_s1_writedata;       // mm_interconnect_0:DDS0_AM_ModPhaseStep_s1_writedata -> DDS0:AM_ModPhaseStep_s1_writedata
	wire         mm_interconnect_0_dds1_am_modphasestep_s1_chipselect;      // mm_interconnect_0:DDS1_AM_ModPhaseStep_s1_chipselect -> DDS1:AM_ModPhaseStep_s1_chipselect
	wire  [31:0] mm_interconnect_0_dds1_am_modphasestep_s1_readdata;        // DDS1:AM_ModPhaseStep_s1_readdata -> mm_interconnect_0:DDS1_AM_ModPhaseStep_s1_readdata
	wire   [1:0] mm_interconnect_0_dds1_am_modphasestep_s1_address;         // mm_interconnect_0:DDS1_AM_ModPhaseStep_s1_address -> DDS1:AM_ModPhaseStep_s1_address
	wire         mm_interconnect_0_dds1_am_modphasestep_s1_write;           // mm_interconnect_0:DDS1_AM_ModPhaseStep_s1_write -> DDS1:AM_ModPhaseStep_s1_write_n
	wire  [31:0] mm_interconnect_0_dds1_am_modphasestep_s1_writedata;       // mm_interconnect_0:DDS1_AM_ModPhaseStep_s1_writedata -> DDS1:AM_ModPhaseStep_s1_writedata
	wire         mm_interconnect_0_lcd_backlight_pwm_s1_chipselect;         // mm_interconnect_0:LCD_BackLight_PWM_s1_chipselect -> LCD:BackLight_PWM_s1_chipselect
	wire  [31:0] mm_interconnect_0_lcd_backlight_pwm_s1_readdata;           // LCD:BackLight_PWM_s1_readdata -> mm_interconnect_0:LCD_BackLight_PWM_s1_readdata
	wire   [1:0] mm_interconnect_0_lcd_backlight_pwm_s1_address;            // mm_interconnect_0:LCD_BackLight_PWM_s1_address -> LCD:BackLight_PWM_s1_address
	wire         mm_interconnect_0_lcd_backlight_pwm_s1_write;              // mm_interconnect_0:LCD_BackLight_PWM_s1_write -> LCD:BackLight_PWM_s1_write_n
	wire  [31:0] mm_interconnect_0_lcd_backlight_pwm_s1_writedata;          // mm_interconnect_0:LCD_BackLight_PWM_s1_writedata -> LCD:BackLight_PWM_s1_writedata
	wire         mm_interconnect_0_lcd_control_s1_chipselect;               // mm_interconnect_0:LCD_Control_s1_chipselect -> LCD:Control_s1_chipselect
	wire  [31:0] mm_interconnect_0_lcd_control_s1_readdata;                 // LCD:Control_s1_readdata -> mm_interconnect_0:LCD_Control_s1_readdata
	wire   [2:0] mm_interconnect_0_lcd_control_s1_address;                  // mm_interconnect_0:LCD_Control_s1_address -> LCD:Control_s1_address
	wire         mm_interconnect_0_lcd_control_s1_write;                    // mm_interconnect_0:LCD_Control_s1_write -> LCD:Control_s1_write_n
	wire  [31:0] mm_interconnect_0_lcd_control_s1_writedata;                // mm_interconnect_0:LCD_Control_s1_writedata -> LCD:Control_s1_writedata
	wire         mm_interconnect_0_lcd_data_s1_chipselect;                  // mm_interconnect_0:LCD_Data_s1_chipselect -> LCD:Data_s1_chipselect
	wire  [31:0] mm_interconnect_0_lcd_data_s1_readdata;                    // LCD:Data_s1_readdata -> mm_interconnect_0:LCD_Data_s1_readdata
	wire   [1:0] mm_interconnect_0_lcd_data_s1_address;                     // mm_interconnect_0:LCD_Data_s1_address -> LCD:Data_s1_address
	wire         mm_interconnect_0_lcd_data_s1_write;                       // mm_interconnect_0:LCD_Data_s1_write -> LCD:Data_s1_write_n
	wire  [31:0] mm_interconnect_0_lcd_data_s1_writedata;                   // mm_interconnect_0:LCD_Data_s1_writedata -> LCD:Data_s1_writedata
	wire         mm_interconnect_0_dds0_fm_moddeviationphase_s1_chipselect; // mm_interconnect_0:DDS0_FM_ModDeviationPhase_s1_chipselect -> DDS0:FM_ModDeviationPhase_s1_chipselect
	wire  [31:0] mm_interconnect_0_dds0_fm_moddeviationphase_s1_readdata;   // DDS0:FM_ModDeviationPhase_s1_readdata -> mm_interconnect_0:DDS0_FM_ModDeviationPhase_s1_readdata
	wire   [1:0] mm_interconnect_0_dds0_fm_moddeviationphase_s1_address;    // mm_interconnect_0:DDS0_FM_ModDeviationPhase_s1_address -> DDS0:FM_ModDeviationPhase_s1_address
	wire         mm_interconnect_0_dds0_fm_moddeviationphase_s1_write;      // mm_interconnect_0:DDS0_FM_ModDeviationPhase_s1_write -> DDS0:FM_ModDeviationPhase_s1_write_n
	wire  [31:0] mm_interconnect_0_dds0_fm_moddeviationphase_s1_writedata;  // mm_interconnect_0:DDS0_FM_ModDeviationPhase_s1_writedata -> DDS0:FM_ModDeviationPhase_s1_writedata
	wire         mm_interconnect_0_dds1_fm_moddeviationphase_s1_chipselect; // mm_interconnect_0:DDS1_FM_ModDeviationPhase_s1_chipselect -> DDS1:FM_ModDeviationPhase_s1_chipselect
	wire  [31:0] mm_interconnect_0_dds1_fm_moddeviationphase_s1_readdata;   // DDS1:FM_ModDeviationPhase_s1_readdata -> mm_interconnect_0:DDS1_FM_ModDeviationPhase_s1_readdata
	wire   [1:0] mm_interconnect_0_dds1_fm_moddeviationphase_s1_address;    // mm_interconnect_0:DDS1_FM_ModDeviationPhase_s1_address -> DDS1:FM_ModDeviationPhase_s1_address
	wire         mm_interconnect_0_dds1_fm_moddeviationphase_s1_write;      // mm_interconnect_0:DDS1_FM_ModDeviationPhase_s1_write -> DDS1:FM_ModDeviationPhase_s1_write_n
	wire  [31:0] mm_interconnect_0_dds1_fm_moddeviationphase_s1_writedata;  // mm_interconnect_0:DDS1_FM_ModDeviationPhase_s1_writedata -> DDS1:FM_ModDeviationPhase_s1_writedata
	wire         mm_interconnect_0_dds0_fm_modphasestep_s1_chipselect;      // mm_interconnect_0:DDS0_FM_ModPhaseStep_s1_chipselect -> DDS0:FM_ModPhaseStep_s1_chipselect
	wire  [31:0] mm_interconnect_0_dds0_fm_modphasestep_s1_readdata;        // DDS0:FM_ModPhaseStep_s1_readdata -> mm_interconnect_0:DDS0_FM_ModPhaseStep_s1_readdata
	wire   [1:0] mm_interconnect_0_dds0_fm_modphasestep_s1_address;         // mm_interconnect_0:DDS0_FM_ModPhaseStep_s1_address -> DDS0:FM_ModPhaseStep_s1_address
	wire         mm_interconnect_0_dds0_fm_modphasestep_s1_write;           // mm_interconnect_0:DDS0_FM_ModPhaseStep_s1_write -> DDS0:FM_ModPhaseStep_s1_write_n
	wire  [31:0] mm_interconnect_0_dds0_fm_modphasestep_s1_writedata;       // mm_interconnect_0:DDS0_FM_ModPhaseStep_s1_writedata -> DDS0:FM_ModPhaseStep_s1_writedata
	wire         mm_interconnect_0_dds1_fm_modphasestep_s1_chipselect;      // mm_interconnect_0:DDS1_FM_ModPhaseStep_s1_chipselect -> DDS1:FM_ModPhaseStep_s1_chipselect
	wire  [31:0] mm_interconnect_0_dds1_fm_modphasestep_s1_readdata;        // DDS1:FM_ModPhaseStep_s1_readdata -> mm_interconnect_0:DDS1_FM_ModPhaseStep_s1_readdata
	wire   [1:0] mm_interconnect_0_dds1_fm_modphasestep_s1_address;         // mm_interconnect_0:DDS1_FM_ModPhaseStep_s1_address -> DDS1:FM_ModPhaseStep_s1_address
	wire         mm_interconnect_0_dds1_fm_modphasestep_s1_write;           // mm_interconnect_0:DDS1_FM_ModPhaseStep_s1_write -> DDS1:FM_ModPhaseStep_s1_write_n
	wire  [31:0] mm_interconnect_0_dds1_fm_modphasestep_s1_writedata;       // mm_interconnect_0:DDS1_FM_ModPhaseStep_s1_writedata -> DDS1:FM_ModPhaseStep_s1_writedata
	wire         mm_interconnect_0_dds0_outputrelay_s1_chipselect;          // mm_interconnect_0:DDS0_OutputRelay_s1_chipselect -> DDS0:OutputRelay_s1_chipselect
	wire  [31:0] mm_interconnect_0_dds0_outputrelay_s1_readdata;            // DDS0:OutputRelay_s1_readdata -> mm_interconnect_0:DDS0_OutputRelay_s1_readdata
	wire   [1:0] mm_interconnect_0_dds0_outputrelay_s1_address;             // mm_interconnect_0:DDS0_OutputRelay_s1_address -> DDS0:OutputRelay_s1_address
	wire         mm_interconnect_0_dds0_outputrelay_s1_write;               // mm_interconnect_0:DDS0_OutputRelay_s1_write -> DDS0:OutputRelay_s1_write_n
	wire  [31:0] mm_interconnect_0_dds0_outputrelay_s1_writedata;           // mm_interconnect_0:DDS0_OutputRelay_s1_writedata -> DDS0:OutputRelay_s1_writedata
	wire         mm_interconnect_0_dds1_outputrelay_s1_chipselect;          // mm_interconnect_0:DDS1_OutputRelay_s1_chipselect -> DDS1:OutputRelay_s1_chipselect
	wire  [31:0] mm_interconnect_0_dds1_outputrelay_s1_readdata;            // DDS1:OutputRelay_s1_readdata -> mm_interconnect_0:DDS1_OutputRelay_s1_readdata
	wire   [1:0] mm_interconnect_0_dds1_outputrelay_s1_address;             // mm_interconnect_0:DDS1_OutputRelay_s1_address -> DDS1:OutputRelay_s1_address
	wire         mm_interconnect_0_dds1_outputrelay_s1_write;               // mm_interconnect_0:DDS1_OutputRelay_s1_write -> DDS1:OutputRelay_s1_write_n
	wire  [31:0] mm_interconnect_0_dds1_outputrelay_s1_writedata;           // mm_interconnect_0:DDS1_OutputRelay_s1_writedata -> DDS1:OutputRelay_s1_writedata
	wire         mm_interconnect_0_dds0_pm_modindex_s1_chipselect;          // mm_interconnect_0:DDS0_PM_ModIndex_s1_chipselect -> DDS0:PM_ModIndex_s1_chipselect
	wire  [31:0] mm_interconnect_0_dds0_pm_modindex_s1_readdata;            // DDS0:PM_ModIndex_s1_readdata -> mm_interconnect_0:DDS0_PM_ModIndex_s1_readdata
	wire   [1:0] mm_interconnect_0_dds0_pm_modindex_s1_address;             // mm_interconnect_0:DDS0_PM_ModIndex_s1_address -> DDS0:PM_ModIndex_s1_address
	wire         mm_interconnect_0_dds0_pm_modindex_s1_write;               // mm_interconnect_0:DDS0_PM_ModIndex_s1_write -> DDS0:PM_ModIndex_s1_write_n
	wire  [31:0] mm_interconnect_0_dds0_pm_modindex_s1_writedata;           // mm_interconnect_0:DDS0_PM_ModIndex_s1_writedata -> DDS0:PM_ModIndex_s1_writedata
	wire         mm_interconnect_0_dds1_pm_modindex_s1_chipselect;          // mm_interconnect_0:DDS1_PM_ModIndex_s1_chipselect -> DDS1:PM_ModIndex_s1_chipselect
	wire  [31:0] mm_interconnect_0_dds1_pm_modindex_s1_readdata;            // DDS1:PM_ModIndex_s1_readdata -> mm_interconnect_0:DDS1_PM_ModIndex_s1_readdata
	wire   [1:0] mm_interconnect_0_dds1_pm_modindex_s1_address;             // mm_interconnect_0:DDS1_PM_ModIndex_s1_address -> DDS1:PM_ModIndex_s1_address
	wire         mm_interconnect_0_dds1_pm_modindex_s1_write;               // mm_interconnect_0:DDS1_PM_ModIndex_s1_write -> DDS1:PM_ModIndex_s1_write_n
	wire  [31:0] mm_interconnect_0_dds1_pm_modindex_s1_writedata;           // mm_interconnect_0:DDS1_PM_ModIndex_s1_writedata -> DDS1:PM_ModIndex_s1_writedata
	wire         mm_interconnect_0_dds0_pm_modphasestep_s1_chipselect;      // mm_interconnect_0:DDS0_PM_ModPhaseStep_s1_chipselect -> DDS0:PM_ModPhaseStep_s1_chipselect
	wire  [31:0] mm_interconnect_0_dds0_pm_modphasestep_s1_readdata;        // DDS0:PM_ModPhaseStep_s1_readdata -> mm_interconnect_0:DDS0_PM_ModPhaseStep_s1_readdata
	wire   [1:0] mm_interconnect_0_dds0_pm_modphasestep_s1_address;         // mm_interconnect_0:DDS0_PM_ModPhaseStep_s1_address -> DDS0:PM_ModPhaseStep_s1_address
	wire         mm_interconnect_0_dds0_pm_modphasestep_s1_write;           // mm_interconnect_0:DDS0_PM_ModPhaseStep_s1_write -> DDS0:PM_ModPhaseStep_s1_write_n
	wire  [31:0] mm_interconnect_0_dds0_pm_modphasestep_s1_writedata;       // mm_interconnect_0:DDS0_PM_ModPhaseStep_s1_writedata -> DDS0:PM_ModPhaseStep_s1_writedata
	wire         mm_interconnect_0_dds1_pm_modphasestep_s1_chipselect;      // mm_interconnect_0:DDS1_PM_ModPhaseStep_s1_chipselect -> DDS1:PM_ModPhaseStep_s1_chipselect
	wire  [31:0] mm_interconnect_0_dds1_pm_modphasestep_s1_readdata;        // DDS1:PM_ModPhaseStep_s1_readdata -> mm_interconnect_0:DDS1_PM_ModPhaseStep_s1_readdata
	wire   [1:0] mm_interconnect_0_dds1_pm_modphasestep_s1_address;         // mm_interconnect_0:DDS1_PM_ModPhaseStep_s1_address -> DDS1:PM_ModPhaseStep_s1_address
	wire         mm_interconnect_0_dds1_pm_modphasestep_s1_write;           // mm_interconnect_0:DDS1_PM_ModPhaseStep_s1_write -> DDS1:PM_ModPhaseStep_s1_write_n
	wire  [31:0] mm_interconnect_0_dds1_pm_modphasestep_s1_writedata;       // mm_interconnect_0:DDS1_PM_ModPhaseStep_s1_writedata -> DDS1:PM_ModPhaseStep_s1_writedata
	wire         mm_interconnect_0_dds0_pwm_amplitude_s1_chipselect;        // mm_interconnect_0:DDS0_PWM_Amplitude_s1_chipselect -> DDS0:PWM_Amplitude_s1_chipselect
	wire  [31:0] mm_interconnect_0_dds0_pwm_amplitude_s1_readdata;          // DDS0:PWM_Amplitude_s1_readdata -> mm_interconnect_0:DDS0_PWM_Amplitude_s1_readdata
	wire   [1:0] mm_interconnect_0_dds0_pwm_amplitude_s1_address;           // mm_interconnect_0:DDS0_PWM_Amplitude_s1_address -> DDS0:PWM_Amplitude_s1_address
	wire         mm_interconnect_0_dds0_pwm_amplitude_s1_write;             // mm_interconnect_0:DDS0_PWM_Amplitude_s1_write -> DDS0:PWM_Amplitude_s1_write_n
	wire  [31:0] mm_interconnect_0_dds0_pwm_amplitude_s1_writedata;         // mm_interconnect_0:DDS0_PWM_Amplitude_s1_writedata -> DDS0:PWM_Amplitude_s1_writedata
	wire         mm_interconnect_0_dds1_pwm_amplitude_s1_chipselect;        // mm_interconnect_0:DDS1_PWM_Amplitude_s1_chipselect -> DDS1:PWM_Amplitude_s1_chipselect
	wire  [31:0] mm_interconnect_0_dds1_pwm_amplitude_s1_readdata;          // DDS1:PWM_Amplitude_s1_readdata -> mm_interconnect_0:DDS1_PWM_Amplitude_s1_readdata
	wire   [1:0] mm_interconnect_0_dds1_pwm_amplitude_s1_address;           // mm_interconnect_0:DDS1_PWM_Amplitude_s1_address -> DDS1:PWM_Amplitude_s1_address
	wire         mm_interconnect_0_dds1_pwm_amplitude_s1_write;             // mm_interconnect_0:DDS1_PWM_Amplitude_s1_write -> DDS1:PWM_Amplitude_s1_write_n
	wire  [31:0] mm_interconnect_0_dds1_pwm_amplitude_s1_writedata;         // mm_interconnect_0:DDS1_PWM_Amplitude_s1_writedata -> DDS1:PWM_Amplitude_s1_writedata
	wire         mm_interconnect_0_dds0_pwm_offset_s1_chipselect;           // mm_interconnect_0:DDS0_PWM_Offset_s1_chipselect -> DDS0:PWM_Offset_s1_chipselect
	wire  [31:0] mm_interconnect_0_dds0_pwm_offset_s1_readdata;             // DDS0:PWM_Offset_s1_readdata -> mm_interconnect_0:DDS0_PWM_Offset_s1_readdata
	wire   [1:0] mm_interconnect_0_dds0_pwm_offset_s1_address;              // mm_interconnect_0:DDS0_PWM_Offset_s1_address -> DDS0:PWM_Offset_s1_address
	wire         mm_interconnect_0_dds0_pwm_offset_s1_write;                // mm_interconnect_0:DDS0_PWM_Offset_s1_write -> DDS0:PWM_Offset_s1_write_n
	wire  [31:0] mm_interconnect_0_dds0_pwm_offset_s1_writedata;            // mm_interconnect_0:DDS0_PWM_Offset_s1_writedata -> DDS0:PWM_Offset_s1_writedata
	wire         mm_interconnect_0_dds1_pwm_offset_s1_chipselect;           // mm_interconnect_0:DDS1_PWM_Offset_s1_chipselect -> DDS1:PWM_Offset_s1_chipselect
	wire  [31:0] mm_interconnect_0_dds1_pwm_offset_s1_readdata;             // DDS1:PWM_Offset_s1_readdata -> mm_interconnect_0:DDS1_PWM_Offset_s1_readdata
	wire   [1:0] mm_interconnect_0_dds1_pwm_offset_s1_address;              // mm_interconnect_0:DDS1_PWM_Offset_s1_address -> DDS1:PWM_Offset_s1_address
	wire         mm_interconnect_0_dds1_pwm_offset_s1_write;                // mm_interconnect_0:DDS1_PWM_Offset_s1_write -> DDS1:PWM_Offset_s1_write_n
	wire  [31:0] mm_interconnect_0_dds1_pwm_offset_s1_writedata;            // mm_interconnect_0:DDS1_PWM_Offset_s1_writedata -> DDS1:PWM_Offset_s1_writedata
	wire         mm_interconnect_0_dds0_phaseoffset_s1_chipselect;          // mm_interconnect_0:DDS0_PhaseOffset_s1_chipselect -> DDS0:PhaseOffset_s1_chipselect
	wire  [31:0] mm_interconnect_0_dds0_phaseoffset_s1_readdata;            // DDS0:PhaseOffset_s1_readdata -> mm_interconnect_0:DDS0_PhaseOffset_s1_readdata
	wire   [1:0] mm_interconnect_0_dds0_phaseoffset_s1_address;             // mm_interconnect_0:DDS0_PhaseOffset_s1_address -> DDS0:PhaseOffset_s1_address
	wire         mm_interconnect_0_dds0_phaseoffset_s1_write;               // mm_interconnect_0:DDS0_PhaseOffset_s1_write -> DDS0:PhaseOffset_s1_write_n
	wire  [31:0] mm_interconnect_0_dds0_phaseoffset_s1_writedata;           // mm_interconnect_0:DDS0_PhaseOffset_s1_writedata -> DDS0:PhaseOffset_s1_writedata
	wire         mm_interconnect_0_dds1_phaseoffset_s1_chipselect;          // mm_interconnect_0:DDS1_PhaseOffset_s1_chipselect -> DDS1:PhaseOffset_s1_chipselect
	wire  [31:0] mm_interconnect_0_dds1_phaseoffset_s1_readdata;            // DDS1:PhaseOffset_s1_readdata -> mm_interconnect_0:DDS1_PhaseOffset_s1_readdata
	wire   [1:0] mm_interconnect_0_dds1_phaseoffset_s1_address;             // mm_interconnect_0:DDS1_PhaseOffset_s1_address -> DDS1:PhaseOffset_s1_address
	wire         mm_interconnect_0_dds1_phaseoffset_s1_write;               // mm_interconnect_0:DDS1_PhaseOffset_s1_write -> DDS1:PhaseOffset_s1_write_n
	wire  [31:0] mm_interconnect_0_dds1_phaseoffset_s1_writedata;           // mm_interconnect_0:DDS1_PhaseOffset_s1_writedata -> DDS1:PhaseOffset_s1_writedata
	wire         mm_interconnect_0_dds0_phasestep_s1_chipselect;            // mm_interconnect_0:DDS0_PhaseStep_s1_chipselect -> DDS0:PhaseStep_s1_chipselect
	wire  [31:0] mm_interconnect_0_dds0_phasestep_s1_readdata;              // DDS0:PhaseStep_s1_readdata -> mm_interconnect_0:DDS0_PhaseStep_s1_readdata
	wire   [1:0] mm_interconnect_0_dds0_phasestep_s1_address;               // mm_interconnect_0:DDS0_PhaseStep_s1_address -> DDS0:PhaseStep_s1_address
	wire         mm_interconnect_0_dds0_phasestep_s1_write;                 // mm_interconnect_0:DDS0_PhaseStep_s1_write -> DDS0:PhaseStep_s1_write_n
	wire  [31:0] mm_interconnect_0_dds0_phasestep_s1_writedata;             // mm_interconnect_0:DDS0_PhaseStep_s1_writedata -> DDS0:PhaseStep_s1_writedata
	wire         mm_interconnect_0_dds1_phasestep_s1_chipselect;            // mm_interconnect_0:DDS1_PhaseStep_s1_chipselect -> DDS1:PhaseStep_s1_chipselect
	wire  [31:0] mm_interconnect_0_dds1_phasestep_s1_readdata;              // DDS1:PhaseStep_s1_readdata -> mm_interconnect_0:DDS1_PhaseStep_s1_readdata
	wire   [1:0] mm_interconnect_0_dds1_phasestep_s1_address;               // mm_interconnect_0:DDS1_PhaseStep_s1_address -> DDS1:PhaseStep_s1_address
	wire         mm_interconnect_0_dds1_phasestep_s1_write;                 // mm_interconnect_0:DDS1_PhaseStep_s1_write -> DDS1:PhaseStep_s1_write_n
	wire  [31:0] mm_interconnect_0_dds1_phasestep_s1_writedata;             // mm_interconnect_0:DDS1_PhaseStep_s1_writedata -> DDS1:PhaseStep_s1_writedata
	wire         mm_interconnect_0_lookup_ram_ram_dds0_am_s1_chipselect;    // mm_interconnect_0:LOOKUP_RAM_RAM_DDS0_AM_s1_chipselect -> LOOKUP_RAM:RAM_DDS0_AM_s1_chipselect
	wire  [15:0] mm_interconnect_0_lookup_ram_ram_dds0_am_s1_readdata;      // LOOKUP_RAM:RAM_DDS0_AM_s1_readdata -> mm_interconnect_0:LOOKUP_RAM_RAM_DDS0_AM_s1_readdata
	wire   [9:0] mm_interconnect_0_lookup_ram_ram_dds0_am_s1_address;       // mm_interconnect_0:LOOKUP_RAM_RAM_DDS0_AM_s1_address -> LOOKUP_RAM:RAM_DDS0_AM_s1_address
	wire   [1:0] mm_interconnect_0_lookup_ram_ram_dds0_am_s1_byteenable;    // mm_interconnect_0:LOOKUP_RAM_RAM_DDS0_AM_s1_byteenable -> LOOKUP_RAM:RAM_DDS0_AM_s1_byteenable
	wire         mm_interconnect_0_lookup_ram_ram_dds0_am_s1_write;         // mm_interconnect_0:LOOKUP_RAM_RAM_DDS0_AM_s1_write -> LOOKUP_RAM:RAM_DDS0_AM_s1_write
	wire  [15:0] mm_interconnect_0_lookup_ram_ram_dds0_am_s1_writedata;     // mm_interconnect_0:LOOKUP_RAM_RAM_DDS0_AM_s1_writedata -> LOOKUP_RAM:RAM_DDS0_AM_s1_writedata
	wire         mm_interconnect_0_lookup_ram_ram_dds0_am_s1_clken;         // mm_interconnect_0:LOOKUP_RAM_RAM_DDS0_AM_s1_clken -> LOOKUP_RAM:RAM_DDS0_AM_s1_clken
	wire         mm_interconnect_0_lookup_ram_ram_dds0_fm_s1_chipselect;    // mm_interconnect_0:LOOKUP_RAM_RAM_DDS0_FM_s1_chipselect -> LOOKUP_RAM:RAM_DDS0_FM_s1_chipselect
	wire  [15:0] mm_interconnect_0_lookup_ram_ram_dds0_fm_s1_readdata;      // LOOKUP_RAM:RAM_DDS0_FM_s1_readdata -> mm_interconnect_0:LOOKUP_RAM_RAM_DDS0_FM_s1_readdata
	wire   [9:0] mm_interconnect_0_lookup_ram_ram_dds0_fm_s1_address;       // mm_interconnect_0:LOOKUP_RAM_RAM_DDS0_FM_s1_address -> LOOKUP_RAM:RAM_DDS0_FM_s1_address
	wire   [1:0] mm_interconnect_0_lookup_ram_ram_dds0_fm_s1_byteenable;    // mm_interconnect_0:LOOKUP_RAM_RAM_DDS0_FM_s1_byteenable -> LOOKUP_RAM:RAM_DDS0_FM_s1_byteenable
	wire         mm_interconnect_0_lookup_ram_ram_dds0_fm_s1_write;         // mm_interconnect_0:LOOKUP_RAM_RAM_DDS0_FM_s1_write -> LOOKUP_RAM:RAM_DDS0_FM_s1_write
	wire  [15:0] mm_interconnect_0_lookup_ram_ram_dds0_fm_s1_writedata;     // mm_interconnect_0:LOOKUP_RAM_RAM_DDS0_FM_s1_writedata -> LOOKUP_RAM:RAM_DDS0_FM_s1_writedata
	wire         mm_interconnect_0_lookup_ram_ram_dds0_fm_s1_clken;         // mm_interconnect_0:LOOKUP_RAM_RAM_DDS0_FM_s1_clken -> LOOKUP_RAM:RAM_DDS0_FM_s1_clken
	wire         mm_interconnect_0_lookup_ram_ram_dds0_s1_chipselect;       // mm_interconnect_0:LOOKUP_RAM_RAM_DDS0_s1_chipselect -> LOOKUP_RAM:RAM_DDS0_s1_chipselect
	wire  [15:0] mm_interconnect_0_lookup_ram_ram_dds0_s1_readdata;         // LOOKUP_RAM:RAM_DDS0_s1_readdata -> mm_interconnect_0:LOOKUP_RAM_RAM_DDS0_s1_readdata
	wire   [9:0] mm_interconnect_0_lookup_ram_ram_dds0_s1_address;          // mm_interconnect_0:LOOKUP_RAM_RAM_DDS0_s1_address -> LOOKUP_RAM:RAM_DDS0_s1_address
	wire   [1:0] mm_interconnect_0_lookup_ram_ram_dds0_s1_byteenable;       // mm_interconnect_0:LOOKUP_RAM_RAM_DDS0_s1_byteenable -> LOOKUP_RAM:RAM_DDS0_s1_byteenable
	wire         mm_interconnect_0_lookup_ram_ram_dds0_s1_write;            // mm_interconnect_0:LOOKUP_RAM_RAM_DDS0_s1_write -> LOOKUP_RAM:RAM_DDS0_s1_write
	wire  [15:0] mm_interconnect_0_lookup_ram_ram_dds0_s1_writedata;        // mm_interconnect_0:LOOKUP_RAM_RAM_DDS0_s1_writedata -> LOOKUP_RAM:RAM_DDS0_s1_writedata
	wire         mm_interconnect_0_lookup_ram_ram_dds0_s1_clken;            // mm_interconnect_0:LOOKUP_RAM_RAM_DDS0_s1_clken -> LOOKUP_RAM:RAM_DDS0_s1_clken
	wire         mm_interconnect_0_lookup_ram_ram_dds1_am_s1_chipselect;    // mm_interconnect_0:LOOKUP_RAM_RAM_DDS1_AM_s1_chipselect -> LOOKUP_RAM:RAM_DDS1_AM_s1_chipselect
	wire  [15:0] mm_interconnect_0_lookup_ram_ram_dds1_am_s1_readdata;      // LOOKUP_RAM:RAM_DDS1_AM_s1_readdata -> mm_interconnect_0:LOOKUP_RAM_RAM_DDS1_AM_s1_readdata
	wire   [9:0] mm_interconnect_0_lookup_ram_ram_dds1_am_s1_address;       // mm_interconnect_0:LOOKUP_RAM_RAM_DDS1_AM_s1_address -> LOOKUP_RAM:RAM_DDS1_AM_s1_address
	wire   [1:0] mm_interconnect_0_lookup_ram_ram_dds1_am_s1_byteenable;    // mm_interconnect_0:LOOKUP_RAM_RAM_DDS1_AM_s1_byteenable -> LOOKUP_RAM:RAM_DDS1_AM_s1_byteenable
	wire         mm_interconnect_0_lookup_ram_ram_dds1_am_s1_write;         // mm_interconnect_0:LOOKUP_RAM_RAM_DDS1_AM_s1_write -> LOOKUP_RAM:RAM_DDS1_AM_s1_write
	wire  [15:0] mm_interconnect_0_lookup_ram_ram_dds1_am_s1_writedata;     // mm_interconnect_0:LOOKUP_RAM_RAM_DDS1_AM_s1_writedata -> LOOKUP_RAM:RAM_DDS1_AM_s1_writedata
	wire         mm_interconnect_0_lookup_ram_ram_dds1_am_s1_clken;         // mm_interconnect_0:LOOKUP_RAM_RAM_DDS1_AM_s1_clken -> LOOKUP_RAM:RAM_DDS1_AM_s1_clken
	wire         mm_interconnect_0_lookup_ram_ram_dds1_fm_s1_chipselect;    // mm_interconnect_0:LOOKUP_RAM_RAM_DDS1_FM_s1_chipselect -> LOOKUP_RAM:RAM_DDS1_FM_s1_chipselect
	wire  [15:0] mm_interconnect_0_lookup_ram_ram_dds1_fm_s1_readdata;      // LOOKUP_RAM:RAM_DDS1_FM_s1_readdata -> mm_interconnect_0:LOOKUP_RAM_RAM_DDS1_FM_s1_readdata
	wire   [9:0] mm_interconnect_0_lookup_ram_ram_dds1_fm_s1_address;       // mm_interconnect_0:LOOKUP_RAM_RAM_DDS1_FM_s1_address -> LOOKUP_RAM:RAM_DDS1_FM_s1_address
	wire   [1:0] mm_interconnect_0_lookup_ram_ram_dds1_fm_s1_byteenable;    // mm_interconnect_0:LOOKUP_RAM_RAM_DDS1_FM_s1_byteenable -> LOOKUP_RAM:RAM_DDS1_FM_s1_byteenable
	wire         mm_interconnect_0_lookup_ram_ram_dds1_fm_s1_write;         // mm_interconnect_0:LOOKUP_RAM_RAM_DDS1_FM_s1_write -> LOOKUP_RAM:RAM_DDS1_FM_s1_write
	wire  [15:0] mm_interconnect_0_lookup_ram_ram_dds1_fm_s1_writedata;     // mm_interconnect_0:LOOKUP_RAM_RAM_DDS1_FM_s1_writedata -> LOOKUP_RAM:RAM_DDS1_FM_s1_writedata
	wire         mm_interconnect_0_lookup_ram_ram_dds1_fm_s1_clken;         // mm_interconnect_0:LOOKUP_RAM_RAM_DDS1_FM_s1_clken -> LOOKUP_RAM:RAM_DDS1_FM_s1_clken
	wire         mm_interconnect_0_lookup_ram_ram_dds1_s1_chipselect;       // mm_interconnect_0:LOOKUP_RAM_RAM_DDS1_s1_chipselect -> LOOKUP_RAM:RAM_DDS1_s1_chipselect
	wire  [15:0] mm_interconnect_0_lookup_ram_ram_dds1_s1_readdata;         // LOOKUP_RAM:RAM_DDS1_s1_readdata -> mm_interconnect_0:LOOKUP_RAM_RAM_DDS1_s1_readdata
	wire   [9:0] mm_interconnect_0_lookup_ram_ram_dds1_s1_address;          // mm_interconnect_0:LOOKUP_RAM_RAM_DDS1_s1_address -> LOOKUP_RAM:RAM_DDS1_s1_address
	wire   [1:0] mm_interconnect_0_lookup_ram_ram_dds1_s1_byteenable;       // mm_interconnect_0:LOOKUP_RAM_RAM_DDS1_s1_byteenable -> LOOKUP_RAM:RAM_DDS1_s1_byteenable
	wire         mm_interconnect_0_lookup_ram_ram_dds1_s1_write;            // mm_interconnect_0:LOOKUP_RAM_RAM_DDS1_s1_write -> LOOKUP_RAM:RAM_DDS1_s1_write
	wire  [15:0] mm_interconnect_0_lookup_ram_ram_dds1_s1_writedata;        // mm_interconnect_0:LOOKUP_RAM_RAM_DDS1_s1_writedata -> LOOKUP_RAM:RAM_DDS1_s1_writedata
	wire         mm_interconnect_0_lookup_ram_ram_dds1_s1_clken;            // mm_interconnect_0:LOOKUP_RAM_RAM_DDS1_s1_clken -> LOOKUP_RAM:RAM_DDS1_s1_clken
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_chipselect -> JTAG_UART:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // JTAG_UART:av_readdata -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // JTAG_UART:av_waitrequest -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_address -> JTAG_UART:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_read -> JTAG_UART:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_write -> JTAG_UART:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_writedata -> JTAG_UART:av_writedata
	wire         mm_interconnect_0_lcd_dma_control_port_slave_chipselect;   // mm_interconnect_0:LCD_DMA_control_port_slave_chipselect -> LCD_DMA:dma_ctl_chipselect
	wire  [14:0] mm_interconnect_0_lcd_dma_control_port_slave_readdata;     // LCD_DMA:dma_ctl_readdata -> mm_interconnect_0:LCD_DMA_control_port_slave_readdata
	wire   [2:0] mm_interconnect_0_lcd_dma_control_port_slave_address;      // mm_interconnect_0:LCD_DMA_control_port_slave_address -> LCD_DMA:dma_ctl_address
	wire         mm_interconnect_0_lcd_dma_control_port_slave_write;        // mm_interconnect_0:LCD_DMA_control_port_slave_write -> LCD_DMA:dma_ctl_write_n
	wire  [14:0] mm_interconnect_0_lcd_dma_control_port_slave_writedata;    // mm_interconnect_0:LCD_DMA_control_port_slave_writedata -> LCD_DMA:dma_ctl_writedata
	wire         mm_interconnect_0_spi_dma_control_port_slave_chipselect;   // mm_interconnect_0:SPI_DMA_control_port_slave_chipselect -> SPI_DMA:dma_ctl_chipselect
	wire  [14:0] mm_interconnect_0_spi_dma_control_port_slave_readdata;     // SPI_DMA:dma_ctl_readdata -> mm_interconnect_0:SPI_DMA_control_port_slave_readdata
	wire   [2:0] mm_interconnect_0_spi_dma_control_port_slave_address;      // mm_interconnect_0:SPI_DMA_control_port_slave_address -> SPI_DMA:dma_ctl_address
	wire         mm_interconnect_0_spi_dma_control_port_slave_write;        // mm_interconnect_0:SPI_DMA_control_port_slave_write -> SPI_DMA:dma_ctl_write_n
	wire  [14:0] mm_interconnect_0_spi_dma_control_port_slave_writedata;    // mm_interconnect_0:SPI_DMA_control_port_slave_writedata -> SPI_DMA:dma_ctl_writedata
	wire  [31:0] mm_interconnect_0_flash_csr_readdata;                      // FLASH:avmm_csr_readdata -> mm_interconnect_0:FLASH_csr_readdata
	wire   [0:0] mm_interconnect_0_flash_csr_address;                       // mm_interconnect_0:FLASH_csr_address -> FLASH:avmm_csr_addr
	wire         mm_interconnect_0_flash_csr_read;                          // mm_interconnect_0:FLASH_csr_read -> FLASH:avmm_csr_read
	wire         mm_interconnect_0_flash_csr_write;                         // mm_interconnect_0:FLASH_csr_write -> FLASH:avmm_csr_write
	wire  [31:0] mm_interconnect_0_flash_csr_writedata;                     // mm_interconnect_0:FLASH_csr_writedata -> FLASH:avmm_csr_writedata
	wire  [31:0] mm_interconnect_0_flash_data_readdata;                     // FLASH:avmm_data_readdata -> mm_interconnect_0:FLASH_data_readdata
	wire         mm_interconnect_0_flash_data_waitrequest;                  // FLASH:avmm_data_waitrequest -> mm_interconnect_0:FLASH_data_waitrequest
	wire  [15:0] mm_interconnect_0_flash_data_address;                      // mm_interconnect_0:FLASH_data_address -> FLASH:avmm_data_addr
	wire         mm_interconnect_0_flash_data_read;                         // mm_interconnect_0:FLASH_data_read -> FLASH:avmm_data_read
	wire         mm_interconnect_0_flash_data_readdatavalid;                // FLASH:avmm_data_readdatavalid -> mm_interconnect_0:FLASH_data_readdatavalid
	wire         mm_interconnect_0_flash_data_write;                        // mm_interconnect_0:FLASH_data_write -> FLASH:avmm_data_write
	wire  [31:0] mm_interconnect_0_flash_data_writedata;                    // mm_interconnect_0:FLASH_data_writedata -> FLASH:avmm_data_writedata
	wire   [3:0] mm_interconnect_0_flash_data_burstcount;                   // mm_interconnect_0:FLASH_data_burstcount -> FLASH:avmm_data_burstcount
	wire  [31:0] mm_interconnect_0_nios_cpu_debug_mem_slave_readdata;       // NIOS_CPU:debug_mem_slave_readdata -> mm_interconnect_0:NIOS_CPU_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios_cpu_debug_mem_slave_waitrequest;    // NIOS_CPU:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOS_CPU_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios_cpu_debug_mem_slave_debugaccess;    // mm_interconnect_0:NIOS_CPU_debug_mem_slave_debugaccess -> NIOS_CPU:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios_cpu_debug_mem_slave_address;        // mm_interconnect_0:NIOS_CPU_debug_mem_slave_address -> NIOS_CPU:debug_mem_slave_address
	wire         mm_interconnect_0_nios_cpu_debug_mem_slave_read;           // mm_interconnect_0:NIOS_CPU_debug_mem_slave_read -> NIOS_CPU:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios_cpu_debug_mem_slave_byteenable;     // mm_interconnect_0:NIOS_CPU_debug_mem_slave_byteenable -> NIOS_CPU:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios_cpu_debug_mem_slave_write;          // mm_interconnect_0:NIOS_CPU_debug_mem_slave_write -> NIOS_CPU:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios_cpu_debug_mem_slave_writedata;      // mm_interconnect_0:NIOS_CPU_debug_mem_slave_writedata -> NIOS_CPU:debug_mem_slave_writedata
	wire         mm_interconnect_0_ram_24k_s1_chipselect;                   // mm_interconnect_0:RAM_24K_s1_chipselect -> RAM_24K:chipselect
	wire  [31:0] mm_interconnect_0_ram_24k_s1_readdata;                     // RAM_24K:readdata -> mm_interconnect_0:RAM_24K_s1_readdata
	wire  [12:0] mm_interconnect_0_ram_24k_s1_address;                      // mm_interconnect_0:RAM_24K_s1_address -> RAM_24K:address
	wire   [3:0] mm_interconnect_0_ram_24k_s1_byteenable;                   // mm_interconnect_0:RAM_24K_s1_byteenable -> RAM_24K:byteenable
	wire         mm_interconnect_0_ram_24k_s1_write;                        // mm_interconnect_0:RAM_24K_s1_write -> RAM_24K:write
	wire  [31:0] mm_interconnect_0_ram_24k_s1_writedata;                    // mm_interconnect_0:RAM_24K_s1_writedata -> RAM_24K:writedata
	wire         mm_interconnect_0_ram_24k_s1_clken;                        // mm_interconnect_0:RAM_24K_s1_clken -> RAM_24K:clken
	wire         mm_interconnect_0_pio_led_debug_s1_chipselect;             // mm_interconnect_0:PIO_LED_DEBUG_s1_chipselect -> PIO_LED_DEBUG:chipselect
	wire  [31:0] mm_interconnect_0_pio_led_debug_s1_readdata;               // PIO_LED_DEBUG:readdata -> mm_interconnect_0:PIO_LED_DEBUG_s1_readdata
	wire   [2:0] mm_interconnect_0_pio_led_debug_s1_address;                // mm_interconnect_0:PIO_LED_DEBUG_s1_address -> PIO_LED_DEBUG:address
	wire         mm_interconnect_0_pio_led_debug_s1_write;                  // mm_interconnect_0:PIO_LED_DEBUG_s1_write -> PIO_LED_DEBUG:write_n
	wire  [31:0] mm_interconnect_0_pio_led_debug_s1_writedata;              // mm_interconnect_0:PIO_LED_DEBUG_s1_writedata -> PIO_LED_DEBUG:writedata
	wire         mm_interconnect_0_timer_delay_32bit_s1_chipselect;         // mm_interconnect_0:TIMER_DELAY_32bit_s1_chipselect -> TIMER_DELAY_32bit:chipselect
	wire  [15:0] mm_interconnect_0_timer_delay_32bit_s1_readdata;           // TIMER_DELAY_32bit:readdata -> mm_interconnect_0:TIMER_DELAY_32bit_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_delay_32bit_s1_address;            // mm_interconnect_0:TIMER_DELAY_32bit_s1_address -> TIMER_DELAY_32bit:address
	wire         mm_interconnect_0_timer_delay_32bit_s1_write;              // mm_interconnect_0:TIMER_DELAY_32bit_s1_write -> TIMER_DELAY_32bit:write_n
	wire  [15:0] mm_interconnect_0_timer_delay_32bit_s1_writedata;          // mm_interconnect_0:TIMER_DELAY_32bit_s1_writedata -> TIMER_DELAY_32bit:writedata
	wire         mm_interconnect_0_keypad_s1_chipselect;                    // mm_interconnect_0:KEYPAD_s1_chipselect -> KEYPAD:chipselect
	wire  [31:0] mm_interconnect_0_keypad_s1_readdata;                      // KEYPAD:readdata -> mm_interconnect_0:KEYPAD_s1_readdata
	wire   [1:0] mm_interconnect_0_keypad_s1_address;                       // mm_interconnect_0:KEYPAD_s1_address -> KEYPAD:address
	wire         mm_interconnect_0_keypad_s1_write;                         // mm_interconnect_0:KEYPAD_s1_write -> KEYPAD:write_n
	wire  [31:0] mm_interconnect_0_keypad_s1_writedata;                     // mm_interconnect_0:KEYPAD_s1_writedata -> KEYPAD:writedata
	wire         mm_interconnect_0_btn_display_s1_chipselect;               // mm_interconnect_0:BTN_DISPLAY_s1_chipselect -> BTN_DISPLAY:chipselect
	wire  [31:0] mm_interconnect_0_btn_display_s1_readdata;                 // BTN_DISPLAY:readdata -> mm_interconnect_0:BTN_DISPLAY_s1_readdata
	wire   [1:0] mm_interconnect_0_btn_display_s1_address;                  // mm_interconnect_0:BTN_DISPLAY_s1_address -> BTN_DISPLAY:address
	wire         mm_interconnect_0_btn_display_s1_write;                    // mm_interconnect_0:BTN_DISPLAY_s1_write -> BTN_DISPLAY:write_n
	wire  [31:0] mm_interconnect_0_btn_display_s1_writedata;                // mm_interconnect_0:BTN_DISPLAY_s1_writedata -> BTN_DISPLAY:writedata
	wire         mm_interconnect_0_btn_encoder_s1_chipselect;               // mm_interconnect_0:BTN_ENCODER_s1_chipselect -> BTN_ENCODER:chipselect
	wire  [31:0] mm_interconnect_0_btn_encoder_s1_readdata;                 // BTN_ENCODER:readdata -> mm_interconnect_0:BTN_ENCODER_s1_readdata
	wire   [1:0] mm_interconnect_0_btn_encoder_s1_address;                  // mm_interconnect_0:BTN_ENCODER_s1_address -> BTN_ENCODER:address
	wire         mm_interconnect_0_btn_encoder_s1_write;                    // mm_interconnect_0:BTN_ENCODER_s1_write -> BTN_ENCODER:write_n
	wire  [31:0] mm_interconnect_0_btn_encoder_s1_writedata;                // mm_interconnect_0:BTN_ENCODER_s1_writedata -> BTN_ENCODER:writedata
	wire         mm_interconnect_0_btn_ch_onoff_s1_chipselect;              // mm_interconnect_0:BTN_CH_ONOFF_s1_chipselect -> BTN_CH_ONOFF:chipselect
	wire  [31:0] mm_interconnect_0_btn_ch_onoff_s1_readdata;                // BTN_CH_ONOFF:readdata -> mm_interconnect_0:BTN_CH_ONOFF_s1_readdata
	wire   [1:0] mm_interconnect_0_btn_ch_onoff_s1_address;                 // mm_interconnect_0:BTN_CH_ONOFF_s1_address -> BTN_CH_ONOFF:address
	wire         mm_interconnect_0_btn_ch_onoff_s1_write;                   // mm_interconnect_0:BTN_CH_ONOFF_s1_write -> BTN_CH_ONOFF:write_n
	wire  [31:0] mm_interconnect_0_btn_ch_onoff_s1_writedata;               // mm_interconnect_0:BTN_CH_ONOFF_s1_writedata -> BTN_CH_ONOFF:writedata
	wire         mm_interconnect_0_dds_reset_s1_chipselect;                 // mm_interconnect_0:DDS_RESET_s1_chipselect -> DDS_RESET:chipselect
	wire  [31:0] mm_interconnect_0_dds_reset_s1_readdata;                   // DDS_RESET:readdata -> mm_interconnect_0:DDS_RESET_s1_readdata
	wire   [1:0] mm_interconnect_0_dds_reset_s1_address;                    // mm_interconnect_0:DDS_RESET_s1_address -> DDS_RESET:address
	wire         mm_interconnect_0_dds_reset_s1_write;                      // mm_interconnect_0:DDS_RESET_s1_write -> DDS_RESET:write_n
	wire  [31:0] mm_interconnect_0_dds_reset_s1_writedata;                  // mm_interconnect_0:DDS_RESET_s1_writedata -> DDS_RESET:writedata
	wire         mm_interconnect_0_lookup_ram_isr_s1_chipselect;            // mm_interconnect_0:LOOKUP_RAM_ISR_s1_chipselect -> LOOKUP_RAM_ISR:chipselect
	wire  [31:0] mm_interconnect_0_lookup_ram_isr_s1_readdata;              // LOOKUP_RAM_ISR:readdata -> mm_interconnect_0:LOOKUP_RAM_ISR_s1_readdata
	wire   [1:0] mm_interconnect_0_lookup_ram_isr_s1_address;               // mm_interconnect_0:LOOKUP_RAM_ISR_s1_address -> LOOKUP_RAM_ISR:address
	wire         mm_interconnect_0_lookup_ram_isr_s1_write;                 // mm_interconnect_0:LOOKUP_RAM_ISR_s1_write -> LOOKUP_RAM_ISR:write_n
	wire  [31:0] mm_interconnect_0_lookup_ram_isr_s1_writedata;             // mm_interconnect_0:LOOKUP_RAM_ISR_s1_writedata -> LOOKUP_RAM_ISR:writedata
	wire         mm_interconnect_0_sd_spi_spi_control_port_chipselect;      // mm_interconnect_0:SD_SPI_spi_control_port_chipselect -> SD_SPI:spi_select
	wire  [15:0] mm_interconnect_0_sd_spi_spi_control_port_readdata;        // SD_SPI:data_to_cpu -> mm_interconnect_0:SD_SPI_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_sd_spi_spi_control_port_address;         // mm_interconnect_0:SD_SPI_spi_control_port_address -> SD_SPI:mem_addr
	wire         mm_interconnect_0_sd_spi_spi_control_port_read;            // mm_interconnect_0:SD_SPI_spi_control_port_read -> SD_SPI:read_n
	wire         mm_interconnect_0_sd_spi_spi_control_port_write;           // mm_interconnect_0:SD_SPI_spi_control_port_write -> SD_SPI:write_n
	wire  [15:0] mm_interconnect_0_sd_spi_spi_control_port_writedata;       // mm_interconnect_0:SD_SPI_spi_control_port_writedata -> SD_SPI:data_from_cpu
	wire         irq_mapper_receiver0_irq;                                  // TIMER_DELAY_32bit:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // KEYPAD:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // BTN_ENCODER:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                  // BTN_DISPLAY:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                  // BTN_CH_ONOFF:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                  // LOOKUP_RAM_ISR:irq -> irq_mapper:receiver5_irq
	wire         irq_mapper_receiver6_irq;                                  // LCD_DMA:dma_ctl_irq -> irq_mapper:receiver6_irq
	wire         irq_mapper_receiver7_irq;                                  // SD_SPI:irq -> irq_mapper:receiver7_irq
	wire         irq_mapper_receiver8_irq;                                  // SPI_DMA:dma_ctl_irq -> irq_mapper:receiver8_irq
	wire         irq_mapper_receiver9_irq;                                  // JTAG_UART:av_irq -> irq_mapper:receiver9_irq
	wire  [31:0] nios_cpu_irq_irq;                                          // irq_mapper:sender_irq -> NIOS_CPU:irq
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [NIOS_CPU:reset_req, RAM_24K:reset_req, rst_translator:reset_req_in]

	NiosII_Processor_BTN_CH_ONOFF btn_ch_onoff (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~cpu_reset),                                   //               reset.reset_n
		.address    (mm_interconnect_0_btn_ch_onoff_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_btn_ch_onoff_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_btn_ch_onoff_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_btn_ch_onoff_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_btn_ch_onoff_s1_readdata),   //                    .readdata
		.in_port    (btn_ch_onoff_export),                          // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                      //                 irq.irq
	);

	NiosII_Processor_BTN_DISPLAY btn_display (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~cpu_reset),                                  //               reset.reset_n
		.address    (mm_interconnect_0_btn_display_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_btn_display_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_btn_display_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_btn_display_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_btn_display_s1_readdata),   //                    .readdata
		.in_port    (btn_display_export),                          // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                     //                 irq.irq
	);

	NiosII_Processor_BTN_ENCODER btn_encoder (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~cpu_reset),                                  //               reset.reset_n
		.address    (mm_interconnect_0_btn_encoder_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_btn_encoder_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_btn_encoder_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_btn_encoder_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_btn_encoder_s1_readdata),   //                    .readdata
		.in_port    (btn_encoder_export),                          // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                     //                 irq.irq
	);

	NiosII_Processor_DDS0 dds0 (
		.AM_ModIndex_clk_clk                             (clk_clk),                                                   //                          AM_ModIndex_clk.clk
		.AM_ModIndex_external_connection_export          (dds0_am_modindex_export),                                   //          AM_ModIndex_external_connection.export
		.AM_ModIndex_reset_reset_n                       (~cpu_reset),                                                //                        AM_ModIndex_reset.reset_n
		.AM_ModIndex_s1_address                          (mm_interconnect_0_dds0_am_modindex_s1_address),             //                           AM_ModIndex_s1.address
		.AM_ModIndex_s1_write_n                          (~mm_interconnect_0_dds0_am_modindex_s1_write),              //                                         .write_n
		.AM_ModIndex_s1_writedata                        (mm_interconnect_0_dds0_am_modindex_s1_writedata),           //                                         .writedata
		.AM_ModIndex_s1_chipselect                       (mm_interconnect_0_dds0_am_modindex_s1_chipselect),          //                                         .chipselect
		.AM_ModIndex_s1_readdata                         (mm_interconnect_0_dds0_am_modindex_s1_readdata),            //                                         .readdata
		.AM_ModPhaseStep_clk_clk                         (clk_clk),                                                   //                      AM_ModPhaseStep_clk.clk
		.AM_ModPhaseStep_external_connection_export      (dds0_am_modphasestep_export),                               //      AM_ModPhaseStep_external_connection.export
		.AM_ModPhaseStep_reset_reset_n                   (~cpu_reset),                                                //                    AM_ModPhaseStep_reset.reset_n
		.AM_ModPhaseStep_s1_address                      (mm_interconnect_0_dds0_am_modphasestep_s1_address),         //                       AM_ModPhaseStep_s1.address
		.AM_ModPhaseStep_s1_write_n                      (~mm_interconnect_0_dds0_am_modphasestep_s1_write),          //                                         .write_n
		.AM_ModPhaseStep_s1_writedata                    (mm_interconnect_0_dds0_am_modphasestep_s1_writedata),       //                                         .writedata
		.AM_ModPhaseStep_s1_chipselect                   (mm_interconnect_0_dds0_am_modphasestep_s1_chipselect),      //                                         .chipselect
		.AM_ModPhaseStep_s1_readdata                     (mm_interconnect_0_dds0_am_modphasestep_s1_readdata),        //                                         .readdata
		.FM_ModDeviationPhase_clk_clk                    (clk_clk),                                                   //                 FM_ModDeviationPhase_clk.clk
		.FM_ModDeviationPhase_external_connection_export (dds0_fm_moddeviationphase_export),                          // FM_ModDeviationPhase_external_connection.export
		.FM_ModDeviationPhase_reset_reset_n              (~cpu_reset),                                                //               FM_ModDeviationPhase_reset.reset_n
		.FM_ModDeviationPhase_s1_address                 (mm_interconnect_0_dds0_fm_moddeviationphase_s1_address),    //                  FM_ModDeviationPhase_s1.address
		.FM_ModDeviationPhase_s1_write_n                 (~mm_interconnect_0_dds0_fm_moddeviationphase_s1_write),     //                                         .write_n
		.FM_ModDeviationPhase_s1_writedata               (mm_interconnect_0_dds0_fm_moddeviationphase_s1_writedata),  //                                         .writedata
		.FM_ModDeviationPhase_s1_chipselect              (mm_interconnect_0_dds0_fm_moddeviationphase_s1_chipselect), //                                         .chipselect
		.FM_ModDeviationPhase_s1_readdata                (mm_interconnect_0_dds0_fm_moddeviationphase_s1_readdata),   //                                         .readdata
		.FM_ModPhaseStep_clk_clk                         (clk_clk),                                                   //                      FM_ModPhaseStep_clk.clk
		.FM_ModPhaseStep_external_connection_export      (dds0_fm_modphasestep_export),                               //      FM_ModPhaseStep_external_connection.export
		.FM_ModPhaseStep_reset_reset_n                   (~cpu_reset),                                                //                    FM_ModPhaseStep_reset.reset_n
		.FM_ModPhaseStep_s1_address                      (mm_interconnect_0_dds0_fm_modphasestep_s1_address),         //                       FM_ModPhaseStep_s1.address
		.FM_ModPhaseStep_s1_write_n                      (~mm_interconnect_0_dds0_fm_modphasestep_s1_write),          //                                         .write_n
		.FM_ModPhaseStep_s1_writedata                    (mm_interconnect_0_dds0_fm_modphasestep_s1_writedata),       //                                         .writedata
		.FM_ModPhaseStep_s1_chipselect                   (mm_interconnect_0_dds0_fm_modphasestep_s1_chipselect),      //                                         .chipselect
		.FM_ModPhaseStep_s1_readdata                     (mm_interconnect_0_dds0_fm_modphasestep_s1_readdata),        //                                         .readdata
		.OutputRelay_clk_clk                             (clk_clk),                                                   //                          OutputRelay_clk.clk
		.OutputRelay_external_connection_export          (dds0_outputrelay_export),                                   //          OutputRelay_external_connection.export
		.OutputRelay_reset_reset_n                       (~cpu_reset),                                                //                        OutputRelay_reset.reset_n
		.OutputRelay_s1_address                          (mm_interconnect_0_dds0_outputrelay_s1_address),             //                           OutputRelay_s1.address
		.OutputRelay_s1_write_n                          (~mm_interconnect_0_dds0_outputrelay_s1_write),              //                                         .write_n
		.OutputRelay_s1_writedata                        (mm_interconnect_0_dds0_outputrelay_s1_writedata),           //                                         .writedata
		.OutputRelay_s1_chipselect                       (mm_interconnect_0_dds0_outputrelay_s1_chipselect),          //                                         .chipselect
		.OutputRelay_s1_readdata                         (mm_interconnect_0_dds0_outputrelay_s1_readdata),            //                                         .readdata
		.PM_ModIndex_clk_clk                             (clk_clk),                                                   //                          PM_ModIndex_clk.clk
		.PM_ModIndex_external_connection_export          (dds0_pm_modindex_export),                                   //          PM_ModIndex_external_connection.export
		.PM_ModIndex_reset_reset_n                       (~cpu_reset),                                                //                        PM_ModIndex_reset.reset_n
		.PM_ModIndex_s1_address                          (mm_interconnect_0_dds0_pm_modindex_s1_address),             //                           PM_ModIndex_s1.address
		.PM_ModIndex_s1_write_n                          (~mm_interconnect_0_dds0_pm_modindex_s1_write),              //                                         .write_n
		.PM_ModIndex_s1_writedata                        (mm_interconnect_0_dds0_pm_modindex_s1_writedata),           //                                         .writedata
		.PM_ModIndex_s1_chipselect                       (mm_interconnect_0_dds0_pm_modindex_s1_chipselect),          //                                         .chipselect
		.PM_ModIndex_s1_readdata                         (mm_interconnect_0_dds0_pm_modindex_s1_readdata),            //                                         .readdata
		.PM_ModPhaseStep_clk_clk                         (clk_clk),                                                   //                      PM_ModPhaseStep_clk.clk
		.PM_ModPhaseStep_external_connection_export      (dds0_pm_modphasestep_export),                               //      PM_ModPhaseStep_external_connection.export
		.PM_ModPhaseStep_reset_reset_n                   (~cpu_reset),                                                //                    PM_ModPhaseStep_reset.reset_n
		.PM_ModPhaseStep_s1_address                      (mm_interconnect_0_dds0_pm_modphasestep_s1_address),         //                       PM_ModPhaseStep_s1.address
		.PM_ModPhaseStep_s1_write_n                      (~mm_interconnect_0_dds0_pm_modphasestep_s1_write),          //                                         .write_n
		.PM_ModPhaseStep_s1_writedata                    (mm_interconnect_0_dds0_pm_modphasestep_s1_writedata),       //                                         .writedata
		.PM_ModPhaseStep_s1_chipselect                   (mm_interconnect_0_dds0_pm_modphasestep_s1_chipselect),      //                                         .chipselect
		.PM_ModPhaseStep_s1_readdata                     (mm_interconnect_0_dds0_pm_modphasestep_s1_readdata),        //                                         .readdata
		.PWM_Amplitude_clk_clk                           (clk_clk),                                                   //                        PWM_Amplitude_clk.clk
		.PWM_Amplitude_external_connection_export        (dds0_pwm_amplitude_export),                                 //        PWM_Amplitude_external_connection.export
		.PWM_Amplitude_reset_reset_n                     (~cpu_reset),                                                //                      PWM_Amplitude_reset.reset_n
		.PWM_Amplitude_s1_address                        (mm_interconnect_0_dds0_pwm_amplitude_s1_address),           //                         PWM_Amplitude_s1.address
		.PWM_Amplitude_s1_write_n                        (~mm_interconnect_0_dds0_pwm_amplitude_s1_write),            //                                         .write_n
		.PWM_Amplitude_s1_writedata                      (mm_interconnect_0_dds0_pwm_amplitude_s1_writedata),         //                                         .writedata
		.PWM_Amplitude_s1_chipselect                     (mm_interconnect_0_dds0_pwm_amplitude_s1_chipselect),        //                                         .chipselect
		.PWM_Amplitude_s1_readdata                       (mm_interconnect_0_dds0_pwm_amplitude_s1_readdata),          //                                         .readdata
		.PWM_Offset_clk_clk                              (clk_clk),                                                   //                           PWM_Offset_clk.clk
		.PWM_Offset_external_connection_export           (dds0_pwm_offset_export),                                    //           PWM_Offset_external_connection.export
		.PWM_Offset_reset_reset_n                        (~cpu_reset),                                                //                         PWM_Offset_reset.reset_n
		.PWM_Offset_s1_address                           (mm_interconnect_0_dds0_pwm_offset_s1_address),              //                            PWM_Offset_s1.address
		.PWM_Offset_s1_write_n                           (~mm_interconnect_0_dds0_pwm_offset_s1_write),               //                                         .write_n
		.PWM_Offset_s1_writedata                         (mm_interconnect_0_dds0_pwm_offset_s1_writedata),            //                                         .writedata
		.PWM_Offset_s1_chipselect                        (mm_interconnect_0_dds0_pwm_offset_s1_chipselect),           //                                         .chipselect
		.PWM_Offset_s1_readdata                          (mm_interconnect_0_dds0_pwm_offset_s1_readdata),             //                                         .readdata
		.PhaseOffset_clk_clk                             (clk_clk),                                                   //                          PhaseOffset_clk.clk
		.PhaseOffset_external_connection_export          (dds0_phaseoffset_export),                                   //          PhaseOffset_external_connection.export
		.PhaseOffset_reset_reset_n                       (~cpu_reset),                                                //                        PhaseOffset_reset.reset_n
		.PhaseOffset_s1_address                          (mm_interconnect_0_dds0_phaseoffset_s1_address),             //                           PhaseOffset_s1.address
		.PhaseOffset_s1_write_n                          (~mm_interconnect_0_dds0_phaseoffset_s1_write),              //                                         .write_n
		.PhaseOffset_s1_writedata                        (mm_interconnect_0_dds0_phaseoffset_s1_writedata),           //                                         .writedata
		.PhaseOffset_s1_chipselect                       (mm_interconnect_0_dds0_phaseoffset_s1_chipselect),          //                                         .chipselect
		.PhaseOffset_s1_readdata                         (mm_interconnect_0_dds0_phaseoffset_s1_readdata),            //                                         .readdata
		.PhaseStep_clk_clk                               (clk_clk),                                                   //                            PhaseStep_clk.clk
		.PhaseStep_external_connection_export            (dds0_phasestep_export),                                     //            PhaseStep_external_connection.export
		.PhaseStep_reset_reset_n                         (~cpu_reset),                                                //                          PhaseStep_reset.reset_n
		.PhaseStep_s1_address                            (mm_interconnect_0_dds0_phasestep_s1_address),               //                             PhaseStep_s1.address
		.PhaseStep_s1_write_n                            (~mm_interconnect_0_dds0_phasestep_s1_write),                //                                         .write_n
		.PhaseStep_s1_writedata                          (mm_interconnect_0_dds0_phasestep_s1_writedata),             //                                         .writedata
		.PhaseStep_s1_chipselect                         (mm_interconnect_0_dds0_phasestep_s1_chipselect),            //                                         .chipselect
		.PhaseStep_s1_readdata                           (mm_interconnect_0_dds0_phasestep_s1_readdata)               //                                         .readdata
	);

	NiosII_Processor_DDS1 dds1 (
		.AM_ModIndex_clk_clk                             (clk_clk),                                                   //                          AM_ModIndex_clk.clk
		.AM_ModIndex_external_connection_export          (dds1_am_modindex_export),                                   //          AM_ModIndex_external_connection.export
		.AM_ModIndex_reset_reset_n                       (~cpu_reset),                                                //                        AM_ModIndex_reset.reset_n
		.AM_ModIndex_s1_address                          (mm_interconnect_0_dds1_am_modindex_s1_address),             //                           AM_ModIndex_s1.address
		.AM_ModIndex_s1_write_n                          (~mm_interconnect_0_dds1_am_modindex_s1_write),              //                                         .write_n
		.AM_ModIndex_s1_writedata                        (mm_interconnect_0_dds1_am_modindex_s1_writedata),           //                                         .writedata
		.AM_ModIndex_s1_chipselect                       (mm_interconnect_0_dds1_am_modindex_s1_chipselect),          //                                         .chipselect
		.AM_ModIndex_s1_readdata                         (mm_interconnect_0_dds1_am_modindex_s1_readdata),            //                                         .readdata
		.AM_ModPhaseStep_clk_clk                         (clk_clk),                                                   //                      AM_ModPhaseStep_clk.clk
		.AM_ModPhaseStep_external_connection_export      (dds1_am_modphasestep_export),                               //      AM_ModPhaseStep_external_connection.export
		.AM_ModPhaseStep_reset_reset_n                   (~cpu_reset),                                                //                    AM_ModPhaseStep_reset.reset_n
		.AM_ModPhaseStep_s1_address                      (mm_interconnect_0_dds1_am_modphasestep_s1_address),         //                       AM_ModPhaseStep_s1.address
		.AM_ModPhaseStep_s1_write_n                      (~mm_interconnect_0_dds1_am_modphasestep_s1_write),          //                                         .write_n
		.AM_ModPhaseStep_s1_writedata                    (mm_interconnect_0_dds1_am_modphasestep_s1_writedata),       //                                         .writedata
		.AM_ModPhaseStep_s1_chipselect                   (mm_interconnect_0_dds1_am_modphasestep_s1_chipselect),      //                                         .chipselect
		.AM_ModPhaseStep_s1_readdata                     (mm_interconnect_0_dds1_am_modphasestep_s1_readdata),        //                                         .readdata
		.FM_ModDeviationPhase_clk_clk                    (clk_clk),                                                   //                 FM_ModDeviationPhase_clk.clk
		.FM_ModDeviationPhase_external_connection_export (dds1_fm_moddeviationphase_export),                          // FM_ModDeviationPhase_external_connection.export
		.FM_ModDeviationPhase_reset_reset_n              (~cpu_reset),                                                //               FM_ModDeviationPhase_reset.reset_n
		.FM_ModDeviationPhase_s1_address                 (mm_interconnect_0_dds1_fm_moddeviationphase_s1_address),    //                  FM_ModDeviationPhase_s1.address
		.FM_ModDeviationPhase_s1_write_n                 (~mm_interconnect_0_dds1_fm_moddeviationphase_s1_write),     //                                         .write_n
		.FM_ModDeviationPhase_s1_writedata               (mm_interconnect_0_dds1_fm_moddeviationphase_s1_writedata),  //                                         .writedata
		.FM_ModDeviationPhase_s1_chipselect              (mm_interconnect_0_dds1_fm_moddeviationphase_s1_chipselect), //                                         .chipselect
		.FM_ModDeviationPhase_s1_readdata                (mm_interconnect_0_dds1_fm_moddeviationphase_s1_readdata),   //                                         .readdata
		.FM_ModPhaseStep_clk_clk                         (clk_clk),                                                   //                      FM_ModPhaseStep_clk.clk
		.FM_ModPhaseStep_external_connection_export      (dds1_fm_modphasestep_export),                               //      FM_ModPhaseStep_external_connection.export
		.FM_ModPhaseStep_reset_reset_n                   (~cpu_reset),                                                //                    FM_ModPhaseStep_reset.reset_n
		.FM_ModPhaseStep_s1_address                      (mm_interconnect_0_dds1_fm_modphasestep_s1_address),         //                       FM_ModPhaseStep_s1.address
		.FM_ModPhaseStep_s1_write_n                      (~mm_interconnect_0_dds1_fm_modphasestep_s1_write),          //                                         .write_n
		.FM_ModPhaseStep_s1_writedata                    (mm_interconnect_0_dds1_fm_modphasestep_s1_writedata),       //                                         .writedata
		.FM_ModPhaseStep_s1_chipselect                   (mm_interconnect_0_dds1_fm_modphasestep_s1_chipselect),      //                                         .chipselect
		.FM_ModPhaseStep_s1_readdata                     (mm_interconnect_0_dds1_fm_modphasestep_s1_readdata),        //                                         .readdata
		.OutputRelay_clk_clk                             (clk_clk),                                                   //                          OutputRelay_clk.clk
		.OutputRelay_external_connection_export          (dds1_outputrelay_export),                                   //          OutputRelay_external_connection.export
		.OutputRelay_reset_reset_n                       (~cpu_reset),                                                //                        OutputRelay_reset.reset_n
		.OutputRelay_s1_address                          (mm_interconnect_0_dds1_outputrelay_s1_address),             //                           OutputRelay_s1.address
		.OutputRelay_s1_write_n                          (~mm_interconnect_0_dds1_outputrelay_s1_write),              //                                         .write_n
		.OutputRelay_s1_writedata                        (mm_interconnect_0_dds1_outputrelay_s1_writedata),           //                                         .writedata
		.OutputRelay_s1_chipselect                       (mm_interconnect_0_dds1_outputrelay_s1_chipselect),          //                                         .chipselect
		.OutputRelay_s1_readdata                         (mm_interconnect_0_dds1_outputrelay_s1_readdata),            //                                         .readdata
		.PM_ModIndex_clk_clk                             (clk_clk),                                                   //                          PM_ModIndex_clk.clk
		.PM_ModIndex_external_connection_export          (dds1_pm_modindex_export),                                   //          PM_ModIndex_external_connection.export
		.PM_ModIndex_reset_reset_n                       (~cpu_reset),                                                //                        PM_ModIndex_reset.reset_n
		.PM_ModIndex_s1_address                          (mm_interconnect_0_dds1_pm_modindex_s1_address),             //                           PM_ModIndex_s1.address
		.PM_ModIndex_s1_write_n                          (~mm_interconnect_0_dds1_pm_modindex_s1_write),              //                                         .write_n
		.PM_ModIndex_s1_writedata                        (mm_interconnect_0_dds1_pm_modindex_s1_writedata),           //                                         .writedata
		.PM_ModIndex_s1_chipselect                       (mm_interconnect_0_dds1_pm_modindex_s1_chipselect),          //                                         .chipselect
		.PM_ModIndex_s1_readdata                         (mm_interconnect_0_dds1_pm_modindex_s1_readdata),            //                                         .readdata
		.PM_ModPhaseStep_clk_clk                         (clk_clk),                                                   //                      PM_ModPhaseStep_clk.clk
		.PM_ModPhaseStep_external_connection_export      (dds1_pm_modphasestep_export),                               //      PM_ModPhaseStep_external_connection.export
		.PM_ModPhaseStep_reset_reset_n                   (~cpu_reset),                                                //                    PM_ModPhaseStep_reset.reset_n
		.PM_ModPhaseStep_s1_address                      (mm_interconnect_0_dds1_pm_modphasestep_s1_address),         //                       PM_ModPhaseStep_s1.address
		.PM_ModPhaseStep_s1_write_n                      (~mm_interconnect_0_dds1_pm_modphasestep_s1_write),          //                                         .write_n
		.PM_ModPhaseStep_s1_writedata                    (mm_interconnect_0_dds1_pm_modphasestep_s1_writedata),       //                                         .writedata
		.PM_ModPhaseStep_s1_chipselect                   (mm_interconnect_0_dds1_pm_modphasestep_s1_chipselect),      //                                         .chipselect
		.PM_ModPhaseStep_s1_readdata                     (mm_interconnect_0_dds1_pm_modphasestep_s1_readdata),        //                                         .readdata
		.PWM_Amplitude_clk_clk                           (clk_clk),                                                   //                        PWM_Amplitude_clk.clk
		.PWM_Amplitude_external_connection_export        (dds1_pwm_amplitude_export),                                 //        PWM_Amplitude_external_connection.export
		.PWM_Amplitude_reset_reset_n                     (~cpu_reset),                                                //                      PWM_Amplitude_reset.reset_n
		.PWM_Amplitude_s1_address                        (mm_interconnect_0_dds1_pwm_amplitude_s1_address),           //                         PWM_Amplitude_s1.address
		.PWM_Amplitude_s1_write_n                        (~mm_interconnect_0_dds1_pwm_amplitude_s1_write),            //                                         .write_n
		.PWM_Amplitude_s1_writedata                      (mm_interconnect_0_dds1_pwm_amplitude_s1_writedata),         //                                         .writedata
		.PWM_Amplitude_s1_chipselect                     (mm_interconnect_0_dds1_pwm_amplitude_s1_chipselect),        //                                         .chipselect
		.PWM_Amplitude_s1_readdata                       (mm_interconnect_0_dds1_pwm_amplitude_s1_readdata),          //                                         .readdata
		.PWM_Offset_clk_clk                              (clk_clk),                                                   //                           PWM_Offset_clk.clk
		.PWM_Offset_external_connection_export           (dds1_pwm_offset_export),                                    //           PWM_Offset_external_connection.export
		.PWM_Offset_reset_reset_n                        (~cpu_reset),                                                //                         PWM_Offset_reset.reset_n
		.PWM_Offset_s1_address                           (mm_interconnect_0_dds1_pwm_offset_s1_address),              //                            PWM_Offset_s1.address
		.PWM_Offset_s1_write_n                           (~mm_interconnect_0_dds1_pwm_offset_s1_write),               //                                         .write_n
		.PWM_Offset_s1_writedata                         (mm_interconnect_0_dds1_pwm_offset_s1_writedata),            //                                         .writedata
		.PWM_Offset_s1_chipselect                        (mm_interconnect_0_dds1_pwm_offset_s1_chipselect),           //                                         .chipselect
		.PWM_Offset_s1_readdata                          (mm_interconnect_0_dds1_pwm_offset_s1_readdata),             //                                         .readdata
		.PhaseOffset_clk_clk                             (clk_clk),                                                   //                          PhaseOffset_clk.clk
		.PhaseOffset_external_connection_export          (dds1_phaseoffset_export),                                   //          PhaseOffset_external_connection.export
		.PhaseOffset_reset_reset_n                       (~cpu_reset),                                                //                        PhaseOffset_reset.reset_n
		.PhaseOffset_s1_address                          (mm_interconnect_0_dds1_phaseoffset_s1_address),             //                           PhaseOffset_s1.address
		.PhaseOffset_s1_write_n                          (~mm_interconnect_0_dds1_phaseoffset_s1_write),              //                                         .write_n
		.PhaseOffset_s1_writedata                        (mm_interconnect_0_dds1_phaseoffset_s1_writedata),           //                                         .writedata
		.PhaseOffset_s1_chipselect                       (mm_interconnect_0_dds1_phaseoffset_s1_chipselect),          //                                         .chipselect
		.PhaseOffset_s1_readdata                         (mm_interconnect_0_dds1_phaseoffset_s1_readdata),            //                                         .readdata
		.PhaseStep_clk_clk                               (clk_clk),                                                   //                            PhaseStep_clk.clk
		.PhaseStep_external_connection_export            (dds1_phasestep_export),                                     //            PhaseStep_external_connection.export
		.PhaseStep_reset_reset_n                         (~cpu_reset),                                                //                          PhaseStep_reset.reset_n
		.PhaseStep_s1_address                            (mm_interconnect_0_dds1_phasestep_s1_address),               //                             PhaseStep_s1.address
		.PhaseStep_s1_write_n                            (~mm_interconnect_0_dds1_phasestep_s1_write),                //                                         .write_n
		.PhaseStep_s1_writedata                          (mm_interconnect_0_dds1_phasestep_s1_writedata),             //                                         .writedata
		.PhaseStep_s1_chipselect                         (mm_interconnect_0_dds1_phasestep_s1_chipselect),            //                                         .chipselect
		.PhaseStep_s1_readdata                           (mm_interconnect_0_dds1_phasestep_s1_readdata)               //                                         .readdata
	);

	NiosII_Processor_DDS_RESET dds_reset (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~cpu_reset),                                //               reset.reset_n
		.address    (mm_interconnect_0_dds_reset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dds_reset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dds_reset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dds_reset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dds_reset_s1_readdata),   //                    .readdata
		.out_port   (dds_reset_export)                           // external_connection.export
	);

	altera_onchip_flash #(
		.INIT_FILENAME                       ("software/DDS_FunctionGen_20Mhz/mem_init/NiosII_Processor_FLASH.hex"),
		.INIT_FILENAME_SIM                   ("software/DDS_FunctionGen_20Mhz/mem_init/hdl_sim/NiosII_Processor_FLASH.dat"),
		.DEVICE_FAMILY                       ("MAX 10"),
		.PART_NAME                           ("10M08SAE144I7G"),
		.DEVICE_ID                           ("08"),
		.SECTOR1_START_ADDR                  (0),
		.SECTOR1_END_ADDR                    (4095),
		.SECTOR2_START_ADDR                  (4096),
		.SECTOR2_END_ADDR                    (8191),
		.SECTOR3_START_ADDR                  (8192),
		.SECTOR3_END_ADDR                    (29183),
		.SECTOR4_START_ADDR                  (29184),
		.SECTOR4_END_ADDR                    (44031),
		.SECTOR5_START_ADDR                  (0),
		.SECTOR5_END_ADDR                    (0),
		.MIN_VALID_ADDR                      (0),
		.MAX_VALID_ADDR                      (44031),
		.MIN_UFM_VALID_ADDR                  (0),
		.MAX_UFM_VALID_ADDR                  (44031),
		.SECTOR1_MAP                         (1),
		.SECTOR2_MAP                         (2),
		.SECTOR3_MAP                         (3),
		.SECTOR4_MAP                         (4),
		.SECTOR5_MAP                         (0),
		.ADDR_RANGE1_END_ADDR                (44031),
		.ADDR_RANGE2_END_ADDR                (44031),
		.ADDR_RANGE1_OFFSET                  (512),
		.ADDR_RANGE2_OFFSET                  (0),
		.ADDR_RANGE3_OFFSET                  (0),
		.AVMM_DATA_ADDR_WIDTH                (16),
		.AVMM_DATA_DATA_WIDTH                (32),
		.AVMM_DATA_BURSTCOUNT_WIDTH          (4),
		.SECTOR_READ_PROTECTION_MODE         (16),
		.FLASH_SEQ_READ_DATA_COUNT           (2),
		.FLASH_ADDR_ALIGNMENT_BITS           (1),
		.FLASH_READ_CYCLE_MAX_INDEX          (4),
		.FLASH_RESET_CYCLE_MAX_INDEX         (25),
		.FLASH_BUSY_TIMEOUT_CYCLE_MAX_INDEX  (120),
		.FLASH_ERASE_TIMEOUT_CYCLE_MAX_INDEX (35000000),
		.FLASH_WRITE_TIMEOUT_CYCLE_MAX_INDEX (30500),
		.PARALLEL_MODE                       (1),
		.READ_AND_WRITE_MODE                 (1),
		.WRAPPING_BURST_MODE                 (0),
		.IS_DUAL_BOOT                        ("False"),
		.IS_ERAM_SKIP                        ("True"),
		.IS_COMPRESSED_IMAGE                 ("True")
	) flash (
		.clock                   (clk_clk),                                    //    clk.clk
		.reset_n                 (~cpu_reset),                                 // nreset.reset_n
		.avmm_data_addr          (mm_interconnect_0_flash_data_address),       //   data.address
		.avmm_data_read          (mm_interconnect_0_flash_data_read),          //       .read
		.avmm_data_writedata     (mm_interconnect_0_flash_data_writedata),     //       .writedata
		.avmm_data_write         (mm_interconnect_0_flash_data_write),         //       .write
		.avmm_data_readdata      (mm_interconnect_0_flash_data_readdata),      //       .readdata
		.avmm_data_waitrequest   (mm_interconnect_0_flash_data_waitrequest),   //       .waitrequest
		.avmm_data_readdatavalid (mm_interconnect_0_flash_data_readdatavalid), //       .readdatavalid
		.avmm_data_burstcount    (mm_interconnect_0_flash_data_burstcount),    //       .burstcount
		.avmm_csr_addr           (mm_interconnect_0_flash_csr_address),        //    csr.address
		.avmm_csr_read           (mm_interconnect_0_flash_csr_read),           //       .read
		.avmm_csr_writedata      (mm_interconnect_0_flash_csr_writedata),      //       .writedata
		.avmm_csr_write          (mm_interconnect_0_flash_csr_write),          //       .write
		.avmm_csr_readdata       (mm_interconnect_0_flash_csr_readdata)        //       .readdata
	);

	NiosII_Processor_JTAG_UART jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~cpu_reset),                                                //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver9_irq)                                   //               irq.irq
	);

	NiosII_Processor_KEYPAD keypad (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~cpu_reset),                             //               reset.reset_n
		.address    (mm_interconnect_0_keypad_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_keypad_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_keypad_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_keypad_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_keypad_s1_readdata),   //                    .readdata
		.in_port    (keypad_input_export),                    // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                //                 irq.irq
	);

	NiosII_Processor_LCD lcd (
		.BackLight_PWM_clk_clk                    (clk_clk),                                           //                 BackLight_PWM_clk.clk
		.BackLight_PWM_external_connection_export (lcd_backlight_pwm_export),                          // BackLight_PWM_external_connection.export
		.BackLight_PWM_reset_reset_n              (~cpu_reset),                                        //               BackLight_PWM_reset.reset_n
		.BackLight_PWM_s1_address                 (mm_interconnect_0_lcd_backlight_pwm_s1_address),    //                  BackLight_PWM_s1.address
		.BackLight_PWM_s1_write_n                 (~mm_interconnect_0_lcd_backlight_pwm_s1_write),     //                                  .write_n
		.BackLight_PWM_s1_writedata               (mm_interconnect_0_lcd_backlight_pwm_s1_writedata),  //                                  .writedata
		.BackLight_PWM_s1_chipselect              (mm_interconnect_0_lcd_backlight_pwm_s1_chipselect), //                                  .chipselect
		.BackLight_PWM_s1_readdata                (mm_interconnect_0_lcd_backlight_pwm_s1_readdata),   //                                  .readdata
		.Control_clk_clk                          (clk_clk),                                           //                       Control_clk.clk
		.Control_external_connection_export       (lcd_control_export),                                //       Control_external_connection.export
		.Control_reset_reset_n                    (~cpu_reset),                                        //                     Control_reset.reset_n
		.Control_s1_address                       (mm_interconnect_0_lcd_control_s1_address),          //                        Control_s1.address
		.Control_s1_write_n                       (~mm_interconnect_0_lcd_control_s1_write),           //                                  .write_n
		.Control_s1_writedata                     (mm_interconnect_0_lcd_control_s1_writedata),        //                                  .writedata
		.Control_s1_chipselect                    (mm_interconnect_0_lcd_control_s1_chipselect),       //                                  .chipselect
		.Control_s1_readdata                      (mm_interconnect_0_lcd_control_s1_readdata),         //                                  .readdata
		.Data_clk_clk                             (clk_clk),                                           //                          Data_clk.clk
		.Data_reset_reset_n                       (~cpu_reset),                                        //                        Data_reset.reset_n
		.Data_s1_address                          (mm_interconnect_0_lcd_data_s1_address),             //                           Data_s1.address
		.Data_s1_write_n                          (~mm_interconnect_0_lcd_data_s1_write),              //                                  .write_n
		.Data_s1_writedata                        (mm_interconnect_0_lcd_data_s1_writedata),           //                                  .writedata
		.Data_s1_chipselect                       (mm_interconnect_0_lcd_data_s1_chipselect),          //                                  .chipselect
		.Data_s1_readdata                         (mm_interconnect_0_lcd_data_s1_readdata),            //                                  .readdata
		.data_external_connection_export          (lcd_data_export)                                    //          data_external_connection.export
	);

	NiosII_Processor_LCD_DMA lcd_dma (
		.clk                (clk_clk),                                                 //                clk.clk
		.system_reset_n     (~cpu_reset),                                              //              reset.reset_n
		.dma_ctl_address    (mm_interconnect_0_lcd_dma_control_port_slave_address),    // control_port_slave.address
		.dma_ctl_chipselect (mm_interconnect_0_lcd_dma_control_port_slave_chipselect), //                   .chipselect
		.dma_ctl_readdata   (mm_interconnect_0_lcd_dma_control_port_slave_readdata),   //                   .readdata
		.dma_ctl_write_n    (~mm_interconnect_0_lcd_dma_control_port_slave_write),     //                   .write_n
		.dma_ctl_writedata  (mm_interconnect_0_lcd_dma_control_port_slave_writedata),  //                   .writedata
		.dma_ctl_irq        (irq_mapper_receiver6_irq),                                //                irq.irq
		.read_address       (lcd_dma_read_master_address),                             //        read_master.address
		.read_chipselect    (lcd_dma_read_master_chipselect),                          //                   .chipselect
		.read_read_n        (lcd_dma_read_master_read),                                //                   .read_n
		.read_readdata      (lcd_dma_read_master_readdata),                            //                   .readdata
		.read_readdatavalid (lcd_dma_read_master_readdatavalid),                       //                   .readdatavalid
		.read_waitrequest   (lcd_dma_read_master_waitrequest),                         //                   .waitrequest
		.write_address      (lcd_dma_address),                                         //       write_master.address
		.write_chipselect   (lcd_dma_chipselect),                                      //                   .chipselect
		.write_waitrequest  (lcd_dma_waitrequest),                                     //                   .waitrequest
		.write_write_n      (lcd_dma_write_n),                                         //                   .write_n
		.write_writedata    (lcd_dma_writedata)                                        //                   .writedata
	);

	NiosII_Processor_LOOKUP_RAM lookup_ram (
		.RAM_DDS0_AM_clk1_clk            (clk_clk),                                                //        RAM_DDS0_AM_clk1.clk
		.RAM_DDS0_AM_reset1_reset        (cpu_reset),                                              //      RAM_DDS0_AM_reset1.reset
		.RAM_DDS0_AM_s1_address          (mm_interconnect_0_lookup_ram_ram_dds0_am_s1_address),    //          RAM_DDS0_AM_s1.address
		.RAM_DDS0_AM_s1_clken            (mm_interconnect_0_lookup_ram_ram_dds0_am_s1_clken),      //                        .clken
		.RAM_DDS0_AM_s1_chipselect       (mm_interconnect_0_lookup_ram_ram_dds0_am_s1_chipselect), //                        .chipselect
		.RAM_DDS0_AM_s1_write            (mm_interconnect_0_lookup_ram_ram_dds0_am_s1_write),      //                        .write
		.RAM_DDS0_AM_s1_readdata         (mm_interconnect_0_lookup_ram_ram_dds0_am_s1_readdata),   //                        .readdata
		.RAM_DDS0_AM_s1_writedata        (mm_interconnect_0_lookup_ram_ram_dds0_am_s1_writedata),  //                        .writedata
		.RAM_DDS0_AM_s1_byteenable       (mm_interconnect_0_lookup_ram_ram_dds0_am_s1_byteenable), //                        .byteenable
		.RAM_DDS0_AM_s2_address          (ram_dds0_am_address),                                    //          RAM_DDS0_AM_s2.address
		.RAM_DDS0_AM_s2_chipselect       (ram_dds0_am_chipselect),                                 //                        .chipselect
		.RAM_DDS0_AM_s2_clken            (ram_dds0_am_clken),                                      //                        .clken
		.RAM_DDS0_AM_s2_write            (ram_dds0_am_write),                                      //                        .write
		.RAM_DDS0_AM_s2_readdata         (ram_dds0_am_readdata),                                   //                        .readdata
		.RAM_DDS0_AM_s2_writedata        (ram_dds0_am_writedata),                                  //                        .writedata
		.RAM_DDS0_AM_s2_byteenable       (ram_dds0_am_byteenable),                                 //                        .byteenable
		.RAM_DDS0_CLK_in_clk_clk         (ram_dds0_clk_clk),                                       //     RAM_DDS0_CLK_in_clk.clk
		.RAM_DDS0_FM_clk1_clk            (clk_clk),                                                //        RAM_DDS0_FM_clk1.clk
		.RAM_DDS0_FM_reset1_reset        (cpu_reset),                                              //      RAM_DDS0_FM_reset1.reset
		.RAM_DDS0_FM_s1_address          (mm_interconnect_0_lookup_ram_ram_dds0_fm_s1_address),    //          RAM_DDS0_FM_s1.address
		.RAM_DDS0_FM_s1_clken            (mm_interconnect_0_lookup_ram_ram_dds0_fm_s1_clken),      //                        .clken
		.RAM_DDS0_FM_s1_chipselect       (mm_interconnect_0_lookup_ram_ram_dds0_fm_s1_chipselect), //                        .chipselect
		.RAM_DDS0_FM_s1_write            (mm_interconnect_0_lookup_ram_ram_dds0_fm_s1_write),      //                        .write
		.RAM_DDS0_FM_s1_readdata         (mm_interconnect_0_lookup_ram_ram_dds0_fm_s1_readdata),   //                        .readdata
		.RAM_DDS0_FM_s1_writedata        (mm_interconnect_0_lookup_ram_ram_dds0_fm_s1_writedata),  //                        .writedata
		.RAM_DDS0_FM_s1_byteenable       (mm_interconnect_0_lookup_ram_ram_dds0_fm_s1_byteenable), //                        .byteenable
		.RAM_DDS0_FM_s2_address          (ram_dds0_fm_address),                                    //          RAM_DDS0_FM_s2.address
		.RAM_DDS0_FM_s2_chipselect       (ram_dds0_fm_chipselect),                                 //                        .chipselect
		.RAM_DDS0_FM_s2_clken            (ram_dds0_fm_clken),                                      //                        .clken
		.RAM_DDS0_FM_s2_write            (ram_dds0_fm_write),                                      //                        .write
		.RAM_DDS0_FM_s2_readdata         (ram_dds0_fm_readdata),                                   //                        .readdata
		.RAM_DDS0_FM_s2_writedata        (ram_dds0_fm_writedata),                                  //                        .writedata
		.RAM_DDS0_FM_s2_byteenable       (ram_dds0_fm_byteenable),                                 //                        .byteenable
		.RAM_DDS0_RESET_in_reset_reset_n (ram_dds0_reset_reset_n),                                 // RAM_DDS0_RESET_in_reset.reset_n
		.RAM_DDS0_clk1_clk               (clk_clk),                                                //           RAM_DDS0_clk1.clk
		.RAM_DDS0_reset1_reset           (cpu_reset),                                              //         RAM_DDS0_reset1.reset
		.RAM_DDS0_s1_address             (mm_interconnect_0_lookup_ram_ram_dds0_s1_address),       //             RAM_DDS0_s1.address
		.RAM_DDS0_s1_clken               (mm_interconnect_0_lookup_ram_ram_dds0_s1_clken),         //                        .clken
		.RAM_DDS0_s1_chipselect          (mm_interconnect_0_lookup_ram_ram_dds0_s1_chipselect),    //                        .chipselect
		.RAM_DDS0_s1_write               (mm_interconnect_0_lookup_ram_ram_dds0_s1_write),         //                        .write
		.RAM_DDS0_s1_readdata            (mm_interconnect_0_lookup_ram_ram_dds0_s1_readdata),      //                        .readdata
		.RAM_DDS0_s1_writedata           (mm_interconnect_0_lookup_ram_ram_dds0_s1_writedata),     //                        .writedata
		.RAM_DDS0_s1_byteenable          (mm_interconnect_0_lookup_ram_ram_dds0_s1_byteenable),    //                        .byteenable
		.RAM_DDS0_s2_address             (ram_dds0_address),                                       //             RAM_DDS0_s2.address
		.RAM_DDS0_s2_chipselect          (ram_dds0_chipselect),                                    //                        .chipselect
		.RAM_DDS0_s2_clken               (ram_dds0_clken),                                         //                        .clken
		.RAM_DDS0_s2_write               (ram_dds0_write),                                         //                        .write
		.RAM_DDS0_s2_readdata            (ram_dds0_readdata),                                      //                        .readdata
		.RAM_DDS0_s2_writedata           (ram_dds0_writedata),                                     //                        .writedata
		.RAM_DDS0_s2_byteenable          (ram_dds0_byteenable),                                    //                        .byteenable
		.RAM_DDS1_AM_clk1_clk            (clk_clk),                                                //        RAM_DDS1_AM_clk1.clk
		.RAM_DDS1_AM_reset1_reset        (cpu_reset),                                              //      RAM_DDS1_AM_reset1.reset
		.RAM_DDS1_AM_s1_address          (mm_interconnect_0_lookup_ram_ram_dds1_am_s1_address),    //          RAM_DDS1_AM_s1.address
		.RAM_DDS1_AM_s1_clken            (mm_interconnect_0_lookup_ram_ram_dds1_am_s1_clken),      //                        .clken
		.RAM_DDS1_AM_s1_chipselect       (mm_interconnect_0_lookup_ram_ram_dds1_am_s1_chipselect), //                        .chipselect
		.RAM_DDS1_AM_s1_write            (mm_interconnect_0_lookup_ram_ram_dds1_am_s1_write),      //                        .write
		.RAM_DDS1_AM_s1_readdata         (mm_interconnect_0_lookup_ram_ram_dds1_am_s1_readdata),   //                        .readdata
		.RAM_DDS1_AM_s1_writedata        (mm_interconnect_0_lookup_ram_ram_dds1_am_s1_writedata),  //                        .writedata
		.RAM_DDS1_AM_s1_byteenable       (mm_interconnect_0_lookup_ram_ram_dds1_am_s1_byteenable), //                        .byteenable
		.RAM_DDS1_AM_s2_address          (ram_dds1_am_address),                                    //          RAM_DDS1_AM_s2.address
		.RAM_DDS1_AM_s2_chipselect       (ram_dds1_am_chipselect),                                 //                        .chipselect
		.RAM_DDS1_AM_s2_clken            (ram_dds1_am_clken),                                      //                        .clken
		.RAM_DDS1_AM_s2_write            (ram_dds1_am_write),                                      //                        .write
		.RAM_DDS1_AM_s2_readdata         (ram_dds1_am_readdata),                                   //                        .readdata
		.RAM_DDS1_AM_s2_writedata        (ram_dds1_am_writedata),                                  //                        .writedata
		.RAM_DDS1_AM_s2_byteenable       (ram_dds1_am_byteenable),                                 //                        .byteenable
		.RAM_DDS1_FM_clk1_clk            (clk_clk),                                                //        RAM_DDS1_FM_clk1.clk
		.RAM_DDS1_FM_reset1_reset        (cpu_reset),                                              //      RAM_DDS1_FM_reset1.reset
		.RAM_DDS1_FM_s1_address          (mm_interconnect_0_lookup_ram_ram_dds1_fm_s1_address),    //          RAM_DDS1_FM_s1.address
		.RAM_DDS1_FM_s1_clken            (mm_interconnect_0_lookup_ram_ram_dds1_fm_s1_clken),      //                        .clken
		.RAM_DDS1_FM_s1_chipselect       (mm_interconnect_0_lookup_ram_ram_dds1_fm_s1_chipselect), //                        .chipselect
		.RAM_DDS1_FM_s1_write            (mm_interconnect_0_lookup_ram_ram_dds1_fm_s1_write),      //                        .write
		.RAM_DDS1_FM_s1_readdata         (mm_interconnect_0_lookup_ram_ram_dds1_fm_s1_readdata),   //                        .readdata
		.RAM_DDS1_FM_s1_writedata        (mm_interconnect_0_lookup_ram_ram_dds1_fm_s1_writedata),  //                        .writedata
		.RAM_DDS1_FM_s1_byteenable       (mm_interconnect_0_lookup_ram_ram_dds1_fm_s1_byteenable), //                        .byteenable
		.RAM_DDS1_FM_s2_address          (ram_dds1_fm_address),                                    //          RAM_DDS1_FM_s2.address
		.RAM_DDS1_FM_s2_chipselect       (ram_dds1_fm_chipselect),                                 //                        .chipselect
		.RAM_DDS1_FM_s2_clken            (ram_dds1_fm_clken),                                      //                        .clken
		.RAM_DDS1_FM_s2_write            (ram_dds1_fm_write),                                      //                        .write
		.RAM_DDS1_FM_s2_readdata         (ram_dds1_fm_readdata),                                   //                        .readdata
		.RAM_DDS1_FM_s2_writedata        (ram_dds1_fm_writedata),                                  //                        .writedata
		.RAM_DDS1_FM_s2_byteenable       (ram_dds1_fm_byteenable),                                 //                        .byteenable
		.RAM_DDS1_clk1_clk               (clk_clk),                                                //           RAM_DDS1_clk1.clk
		.RAM_DDS1_reset1_reset           (cpu_reset),                                              //         RAM_DDS1_reset1.reset
		.RAM_DDS1_s1_address             (mm_interconnect_0_lookup_ram_ram_dds1_s1_address),       //             RAM_DDS1_s1.address
		.RAM_DDS1_s1_clken               (mm_interconnect_0_lookup_ram_ram_dds1_s1_clken),         //                        .clken
		.RAM_DDS1_s1_chipselect          (mm_interconnect_0_lookup_ram_ram_dds1_s1_chipselect),    //                        .chipselect
		.RAM_DDS1_s1_write               (mm_interconnect_0_lookup_ram_ram_dds1_s1_write),         //                        .write
		.RAM_DDS1_s1_readdata            (mm_interconnect_0_lookup_ram_ram_dds1_s1_readdata),      //                        .readdata
		.RAM_DDS1_s1_writedata           (mm_interconnect_0_lookup_ram_ram_dds1_s1_writedata),     //                        .writedata
		.RAM_DDS1_s1_byteenable          (mm_interconnect_0_lookup_ram_ram_dds1_s1_byteenable),    //                        .byteenable
		.RAM_DDS1_s2_address             (ram_dds1_address),                                       //             RAM_DDS1_s2.address
		.RAM_DDS1_s2_chipselect          (ram_dds1_chipselect),                                    //                        .chipselect
		.RAM_DDS1_s2_clken               (ram_dds1_clken),                                         //                        .clken
		.RAM_DDS1_s2_write               (ram_dds1_write),                                         //                        .write
		.RAM_DDS1_s2_readdata            (ram_dds1_readdata),                                      //                        .readdata
		.RAM_DDS1_s2_writedata           (ram_dds1_writedata),                                     //                        .writedata
		.RAM_DDS1_s2_byteenable          (ram_dds1_byteenable)                                     //                        .byteenable
	);

	NiosII_Processor_LOOKUP_RAM_ISR lookup_ram_isr (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~cpu_reset),                                     //               reset.reset_n
		.address    (mm_interconnect_0_lookup_ram_isr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lookup_ram_isr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lookup_ram_isr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lookup_ram_isr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lookup_ram_isr_s1_readdata),   //                    .readdata
		.in_port    (lookup_ram_isr_1_export),                        // external_connection.export
		.irq        (irq_mapper_receiver5_irq)                        //                 irq.irq
	);

	NiosII_Processor_NIOS_CPU nios_cpu (
		.clk                                 (clk_clk),                                                //                       clk.clk
		.reset_n                             (~cpu_reset),                                             //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios_cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios_cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios_cpu_data_master_read),                              //                          .read
		.d_readdata                          (nios_cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios_cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios_cpu_data_master_write),                             //                          .write
		.d_writedata                         (nios_cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios_cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios_cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios_cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (nios_cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios_cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios_cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios_cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                        // custom_instruction_master.readra
	);

	NiosII_Processor_PIO_LED_DEBUG pio_led_debug (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~cpu_reset),                                    //               reset.reset_n
		.address    (mm_interconnect_0_pio_led_debug_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_led_debug_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_led_debug_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_led_debug_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_led_debug_s1_readdata),   //                    .readdata
		.out_port   (led_debug_export)                               // external_connection.export
	);

	NiosII_Processor_RAM_24K ram_24k (
		.clk        (clk_clk),                                 //   clk1.clk
		.address    (mm_interconnect_0_ram_24k_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_24k_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_24k_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_24k_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_24k_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_24k_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_24k_s1_byteenable), //       .byteenable
		.reset      (cpu_reset),                               // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),      //       .reset_req
		.freeze     (1'b0)                                     // (terminated)
	);

	NiosII_Processor_SD_SPI sd_spi (
		.clk           (clk_clk),                                              //              clk.clk
		.reset_n       (~cpu_reset),                                           //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_sd_spi_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_sd_spi_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_sd_spi_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_sd_spi_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_sd_spi_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_sd_spi_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver7_irq),                             //              irq.irq
		.MISO          (sd_spi_MISO),                                          //         external.export
		.MOSI          (sd_spi_MOSI),                                          //                 .export
		.SCLK          (sd_spi_SCLK),                                          //                 .export
		.SS_n          (sd_spi_SS_n)                                           //                 .export
	);

	NiosII_Processor_SPI_DMA spi_dma (
		.clk                (clk_clk),                                                 //                clk.clk
		.system_reset_n     (~cpu_reset),                                              //              reset.reset_n
		.dma_ctl_address    (mm_interconnect_0_spi_dma_control_port_slave_address),    // control_port_slave.address
		.dma_ctl_chipselect (mm_interconnect_0_spi_dma_control_port_slave_chipselect), //                   .chipselect
		.dma_ctl_readdata   (mm_interconnect_0_spi_dma_control_port_slave_readdata),   //                   .readdata
		.dma_ctl_write_n    (~mm_interconnect_0_spi_dma_control_port_slave_write),     //                   .write_n
		.dma_ctl_writedata  (mm_interconnect_0_spi_dma_control_port_slave_writedata),  //                   .writedata
		.dma_ctl_irq        (irq_mapper_receiver8_irq),                                //                irq.irq
		.read_address       (spi_dma_address),                                         //        read_master.address
		.read_chipselect    (spi_dma_chipselect),                                      //                   .chipselect
		.read_read_n        (spi_dma_read_n),                                          //                   .read_n
		.read_readdata      (spi_dma_readdata),                                        //                   .readdata
		.read_readdatavalid (spi_dma_readdatavalid),                                   //                   .readdatavalid
		.read_waitrequest   (spi_dma_waitrequest),                                     //                   .waitrequest
		.write_address      (spi_dma_write_master_address),                            //       write_master.address
		.write_chipselect   (spi_dma_write_master_chipselect),                         //                   .chipselect
		.write_waitrequest  (spi_dma_write_master_waitrequest),                        //                   .waitrequest
		.write_write_n      (spi_dma_write_master_write),                              //                   .write_n
		.write_writedata    (spi_dma_write_master_writedata)                           //                   .writedata
	);

	NiosII_Processor_TIMER_DELAY_32bit timer_delay_32bit (
		.clk        (clk_clk),                                           //   clk.clk
		.reset_n    (~cpu_reset),                                        // reset.reset_n
		.address    (mm_interconnect_0_timer_delay_32bit_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_delay_32bit_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_delay_32bit_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_delay_32bit_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_delay_32bit_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                           //   irq.irq
	);

	NiosII_Processor_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                              (clk_clk),                                                   //                            clk_0_clk.clk
		.NIOS_CPU_reset_reset_bridge_in_reset_reset (cpu_reset),                                                 // NIOS_CPU_reset_reset_bridge_in_reset.reset
		.LCD_DMA_read_master_address                (lcd_dma_read_master_address),                               //                  LCD_DMA_read_master.address
		.LCD_DMA_read_master_waitrequest            (lcd_dma_read_master_waitrequest),                           //                                     .waitrequest
		.LCD_DMA_read_master_chipselect             (lcd_dma_read_master_chipselect),                            //                                     .chipselect
		.LCD_DMA_read_master_read                   (~lcd_dma_read_master_read),                                 //                                     .read
		.LCD_DMA_read_master_readdata               (lcd_dma_read_master_readdata),                              //                                     .readdata
		.LCD_DMA_read_master_readdatavalid          (lcd_dma_read_master_readdatavalid),                         //                                     .readdatavalid
		.NIOS_CPU_data_master_address               (nios_cpu_data_master_address),                              //                 NIOS_CPU_data_master.address
		.NIOS_CPU_data_master_waitrequest           (nios_cpu_data_master_waitrequest),                          //                                     .waitrequest
		.NIOS_CPU_data_master_byteenable            (nios_cpu_data_master_byteenable),                           //                                     .byteenable
		.NIOS_CPU_data_master_read                  (nios_cpu_data_master_read),                                 //                                     .read
		.NIOS_CPU_data_master_readdata              (nios_cpu_data_master_readdata),                             //                                     .readdata
		.NIOS_CPU_data_master_write                 (nios_cpu_data_master_write),                                //                                     .write
		.NIOS_CPU_data_master_writedata             (nios_cpu_data_master_writedata),                            //                                     .writedata
		.NIOS_CPU_data_master_debugaccess           (nios_cpu_data_master_debugaccess),                          //                                     .debugaccess
		.NIOS_CPU_instruction_master_address        (nios_cpu_instruction_master_address),                       //          NIOS_CPU_instruction_master.address
		.NIOS_CPU_instruction_master_waitrequest    (nios_cpu_instruction_master_waitrequest),                   //                                     .waitrequest
		.NIOS_CPU_instruction_master_read           (nios_cpu_instruction_master_read),                          //                                     .read
		.NIOS_CPU_instruction_master_readdata       (nios_cpu_instruction_master_readdata),                      //                                     .readdata
		.SPI_DMA_write_master_address               (spi_dma_write_master_address),                              //                 SPI_DMA_write_master.address
		.SPI_DMA_write_master_waitrequest           (spi_dma_write_master_waitrequest),                          //                                     .waitrequest
		.SPI_DMA_write_master_chipselect            (spi_dma_write_master_chipselect),                           //                                     .chipselect
		.SPI_DMA_write_master_write                 (~spi_dma_write_master_write),                               //                                     .write
		.SPI_DMA_write_master_writedata             (spi_dma_write_master_writedata),                            //                                     .writedata
		.BTN_CH_ONOFF_s1_address                    (mm_interconnect_0_btn_ch_onoff_s1_address),                 //                      BTN_CH_ONOFF_s1.address
		.BTN_CH_ONOFF_s1_write                      (mm_interconnect_0_btn_ch_onoff_s1_write),                   //                                     .write
		.BTN_CH_ONOFF_s1_readdata                   (mm_interconnect_0_btn_ch_onoff_s1_readdata),                //                                     .readdata
		.BTN_CH_ONOFF_s1_writedata                  (mm_interconnect_0_btn_ch_onoff_s1_writedata),               //                                     .writedata
		.BTN_CH_ONOFF_s1_chipselect                 (mm_interconnect_0_btn_ch_onoff_s1_chipselect),              //                                     .chipselect
		.BTN_DISPLAY_s1_address                     (mm_interconnect_0_btn_display_s1_address),                  //                       BTN_DISPLAY_s1.address
		.BTN_DISPLAY_s1_write                       (mm_interconnect_0_btn_display_s1_write),                    //                                     .write
		.BTN_DISPLAY_s1_readdata                    (mm_interconnect_0_btn_display_s1_readdata),                 //                                     .readdata
		.BTN_DISPLAY_s1_writedata                   (mm_interconnect_0_btn_display_s1_writedata),                //                                     .writedata
		.BTN_DISPLAY_s1_chipselect                  (mm_interconnect_0_btn_display_s1_chipselect),               //                                     .chipselect
		.BTN_ENCODER_s1_address                     (mm_interconnect_0_btn_encoder_s1_address),                  //                       BTN_ENCODER_s1.address
		.BTN_ENCODER_s1_write                       (mm_interconnect_0_btn_encoder_s1_write),                    //                                     .write
		.BTN_ENCODER_s1_readdata                    (mm_interconnect_0_btn_encoder_s1_readdata),                 //                                     .readdata
		.BTN_ENCODER_s1_writedata                   (mm_interconnect_0_btn_encoder_s1_writedata),                //                                     .writedata
		.BTN_ENCODER_s1_chipselect                  (mm_interconnect_0_btn_encoder_s1_chipselect),               //                                     .chipselect
		.DDS0_AM_ModIndex_s1_address                (mm_interconnect_0_dds0_am_modindex_s1_address),             //                  DDS0_AM_ModIndex_s1.address
		.DDS0_AM_ModIndex_s1_write                  (mm_interconnect_0_dds0_am_modindex_s1_write),               //                                     .write
		.DDS0_AM_ModIndex_s1_readdata               (mm_interconnect_0_dds0_am_modindex_s1_readdata),            //                                     .readdata
		.DDS0_AM_ModIndex_s1_writedata              (mm_interconnect_0_dds0_am_modindex_s1_writedata),           //                                     .writedata
		.DDS0_AM_ModIndex_s1_chipselect             (mm_interconnect_0_dds0_am_modindex_s1_chipselect),          //                                     .chipselect
		.DDS0_AM_ModPhaseStep_s1_address            (mm_interconnect_0_dds0_am_modphasestep_s1_address),         //              DDS0_AM_ModPhaseStep_s1.address
		.DDS0_AM_ModPhaseStep_s1_write              (mm_interconnect_0_dds0_am_modphasestep_s1_write),           //                                     .write
		.DDS0_AM_ModPhaseStep_s1_readdata           (mm_interconnect_0_dds0_am_modphasestep_s1_readdata),        //                                     .readdata
		.DDS0_AM_ModPhaseStep_s1_writedata          (mm_interconnect_0_dds0_am_modphasestep_s1_writedata),       //                                     .writedata
		.DDS0_AM_ModPhaseStep_s1_chipselect         (mm_interconnect_0_dds0_am_modphasestep_s1_chipselect),      //                                     .chipselect
		.DDS0_FM_ModDeviationPhase_s1_address       (mm_interconnect_0_dds0_fm_moddeviationphase_s1_address),    //         DDS0_FM_ModDeviationPhase_s1.address
		.DDS0_FM_ModDeviationPhase_s1_write         (mm_interconnect_0_dds0_fm_moddeviationphase_s1_write),      //                                     .write
		.DDS0_FM_ModDeviationPhase_s1_readdata      (mm_interconnect_0_dds0_fm_moddeviationphase_s1_readdata),   //                                     .readdata
		.DDS0_FM_ModDeviationPhase_s1_writedata     (mm_interconnect_0_dds0_fm_moddeviationphase_s1_writedata),  //                                     .writedata
		.DDS0_FM_ModDeviationPhase_s1_chipselect    (mm_interconnect_0_dds0_fm_moddeviationphase_s1_chipselect), //                                     .chipselect
		.DDS0_FM_ModPhaseStep_s1_address            (mm_interconnect_0_dds0_fm_modphasestep_s1_address),         //              DDS0_FM_ModPhaseStep_s1.address
		.DDS0_FM_ModPhaseStep_s1_write              (mm_interconnect_0_dds0_fm_modphasestep_s1_write),           //                                     .write
		.DDS0_FM_ModPhaseStep_s1_readdata           (mm_interconnect_0_dds0_fm_modphasestep_s1_readdata),        //                                     .readdata
		.DDS0_FM_ModPhaseStep_s1_writedata          (mm_interconnect_0_dds0_fm_modphasestep_s1_writedata),       //                                     .writedata
		.DDS0_FM_ModPhaseStep_s1_chipselect         (mm_interconnect_0_dds0_fm_modphasestep_s1_chipselect),      //                                     .chipselect
		.DDS0_OutputRelay_s1_address                (mm_interconnect_0_dds0_outputrelay_s1_address),             //                  DDS0_OutputRelay_s1.address
		.DDS0_OutputRelay_s1_write                  (mm_interconnect_0_dds0_outputrelay_s1_write),               //                                     .write
		.DDS0_OutputRelay_s1_readdata               (mm_interconnect_0_dds0_outputrelay_s1_readdata),            //                                     .readdata
		.DDS0_OutputRelay_s1_writedata              (mm_interconnect_0_dds0_outputrelay_s1_writedata),           //                                     .writedata
		.DDS0_OutputRelay_s1_chipselect             (mm_interconnect_0_dds0_outputrelay_s1_chipselect),          //                                     .chipselect
		.DDS0_PhaseOffset_s1_address                (mm_interconnect_0_dds0_phaseoffset_s1_address),             //                  DDS0_PhaseOffset_s1.address
		.DDS0_PhaseOffset_s1_write                  (mm_interconnect_0_dds0_phaseoffset_s1_write),               //                                     .write
		.DDS0_PhaseOffset_s1_readdata               (mm_interconnect_0_dds0_phaseoffset_s1_readdata),            //                                     .readdata
		.DDS0_PhaseOffset_s1_writedata              (mm_interconnect_0_dds0_phaseoffset_s1_writedata),           //                                     .writedata
		.DDS0_PhaseOffset_s1_chipselect             (mm_interconnect_0_dds0_phaseoffset_s1_chipselect),          //                                     .chipselect
		.DDS0_PhaseStep_s1_address                  (mm_interconnect_0_dds0_phasestep_s1_address),               //                    DDS0_PhaseStep_s1.address
		.DDS0_PhaseStep_s1_write                    (mm_interconnect_0_dds0_phasestep_s1_write),                 //                                     .write
		.DDS0_PhaseStep_s1_readdata                 (mm_interconnect_0_dds0_phasestep_s1_readdata),              //                                     .readdata
		.DDS0_PhaseStep_s1_writedata                (mm_interconnect_0_dds0_phasestep_s1_writedata),             //                                     .writedata
		.DDS0_PhaseStep_s1_chipselect               (mm_interconnect_0_dds0_phasestep_s1_chipselect),            //                                     .chipselect
		.DDS0_PM_ModIndex_s1_address                (mm_interconnect_0_dds0_pm_modindex_s1_address),             //                  DDS0_PM_ModIndex_s1.address
		.DDS0_PM_ModIndex_s1_write                  (mm_interconnect_0_dds0_pm_modindex_s1_write),               //                                     .write
		.DDS0_PM_ModIndex_s1_readdata               (mm_interconnect_0_dds0_pm_modindex_s1_readdata),            //                                     .readdata
		.DDS0_PM_ModIndex_s1_writedata              (mm_interconnect_0_dds0_pm_modindex_s1_writedata),           //                                     .writedata
		.DDS0_PM_ModIndex_s1_chipselect             (mm_interconnect_0_dds0_pm_modindex_s1_chipselect),          //                                     .chipselect
		.DDS0_PM_ModPhaseStep_s1_address            (mm_interconnect_0_dds0_pm_modphasestep_s1_address),         //              DDS0_PM_ModPhaseStep_s1.address
		.DDS0_PM_ModPhaseStep_s1_write              (mm_interconnect_0_dds0_pm_modphasestep_s1_write),           //                                     .write
		.DDS0_PM_ModPhaseStep_s1_readdata           (mm_interconnect_0_dds0_pm_modphasestep_s1_readdata),        //                                     .readdata
		.DDS0_PM_ModPhaseStep_s1_writedata          (mm_interconnect_0_dds0_pm_modphasestep_s1_writedata),       //                                     .writedata
		.DDS0_PM_ModPhaseStep_s1_chipselect         (mm_interconnect_0_dds0_pm_modphasestep_s1_chipselect),      //                                     .chipselect
		.DDS0_PWM_Amplitude_s1_address              (mm_interconnect_0_dds0_pwm_amplitude_s1_address),           //                DDS0_PWM_Amplitude_s1.address
		.DDS0_PWM_Amplitude_s1_write                (mm_interconnect_0_dds0_pwm_amplitude_s1_write),             //                                     .write
		.DDS0_PWM_Amplitude_s1_readdata             (mm_interconnect_0_dds0_pwm_amplitude_s1_readdata),          //                                     .readdata
		.DDS0_PWM_Amplitude_s1_writedata            (mm_interconnect_0_dds0_pwm_amplitude_s1_writedata),         //                                     .writedata
		.DDS0_PWM_Amplitude_s1_chipselect           (mm_interconnect_0_dds0_pwm_amplitude_s1_chipselect),        //                                     .chipselect
		.DDS0_PWM_Offset_s1_address                 (mm_interconnect_0_dds0_pwm_offset_s1_address),              //                   DDS0_PWM_Offset_s1.address
		.DDS0_PWM_Offset_s1_write                   (mm_interconnect_0_dds0_pwm_offset_s1_write),                //                                     .write
		.DDS0_PWM_Offset_s1_readdata                (mm_interconnect_0_dds0_pwm_offset_s1_readdata),             //                                     .readdata
		.DDS0_PWM_Offset_s1_writedata               (mm_interconnect_0_dds0_pwm_offset_s1_writedata),            //                                     .writedata
		.DDS0_PWM_Offset_s1_chipselect              (mm_interconnect_0_dds0_pwm_offset_s1_chipselect),           //                                     .chipselect
		.DDS1_AM_ModIndex_s1_address                (mm_interconnect_0_dds1_am_modindex_s1_address),             //                  DDS1_AM_ModIndex_s1.address
		.DDS1_AM_ModIndex_s1_write                  (mm_interconnect_0_dds1_am_modindex_s1_write),               //                                     .write
		.DDS1_AM_ModIndex_s1_readdata               (mm_interconnect_0_dds1_am_modindex_s1_readdata),            //                                     .readdata
		.DDS1_AM_ModIndex_s1_writedata              (mm_interconnect_0_dds1_am_modindex_s1_writedata),           //                                     .writedata
		.DDS1_AM_ModIndex_s1_chipselect             (mm_interconnect_0_dds1_am_modindex_s1_chipselect),          //                                     .chipselect
		.DDS1_AM_ModPhaseStep_s1_address            (mm_interconnect_0_dds1_am_modphasestep_s1_address),         //              DDS1_AM_ModPhaseStep_s1.address
		.DDS1_AM_ModPhaseStep_s1_write              (mm_interconnect_0_dds1_am_modphasestep_s1_write),           //                                     .write
		.DDS1_AM_ModPhaseStep_s1_readdata           (mm_interconnect_0_dds1_am_modphasestep_s1_readdata),        //                                     .readdata
		.DDS1_AM_ModPhaseStep_s1_writedata          (mm_interconnect_0_dds1_am_modphasestep_s1_writedata),       //                                     .writedata
		.DDS1_AM_ModPhaseStep_s1_chipselect         (mm_interconnect_0_dds1_am_modphasestep_s1_chipselect),      //                                     .chipselect
		.DDS1_FM_ModDeviationPhase_s1_address       (mm_interconnect_0_dds1_fm_moddeviationphase_s1_address),    //         DDS1_FM_ModDeviationPhase_s1.address
		.DDS1_FM_ModDeviationPhase_s1_write         (mm_interconnect_0_dds1_fm_moddeviationphase_s1_write),      //                                     .write
		.DDS1_FM_ModDeviationPhase_s1_readdata      (mm_interconnect_0_dds1_fm_moddeviationphase_s1_readdata),   //                                     .readdata
		.DDS1_FM_ModDeviationPhase_s1_writedata     (mm_interconnect_0_dds1_fm_moddeviationphase_s1_writedata),  //                                     .writedata
		.DDS1_FM_ModDeviationPhase_s1_chipselect    (mm_interconnect_0_dds1_fm_moddeviationphase_s1_chipselect), //                                     .chipselect
		.DDS1_FM_ModPhaseStep_s1_address            (mm_interconnect_0_dds1_fm_modphasestep_s1_address),         //              DDS1_FM_ModPhaseStep_s1.address
		.DDS1_FM_ModPhaseStep_s1_write              (mm_interconnect_0_dds1_fm_modphasestep_s1_write),           //                                     .write
		.DDS1_FM_ModPhaseStep_s1_readdata           (mm_interconnect_0_dds1_fm_modphasestep_s1_readdata),        //                                     .readdata
		.DDS1_FM_ModPhaseStep_s1_writedata          (mm_interconnect_0_dds1_fm_modphasestep_s1_writedata),       //                                     .writedata
		.DDS1_FM_ModPhaseStep_s1_chipselect         (mm_interconnect_0_dds1_fm_modphasestep_s1_chipselect),      //                                     .chipselect
		.DDS1_OutputRelay_s1_address                (mm_interconnect_0_dds1_outputrelay_s1_address),             //                  DDS1_OutputRelay_s1.address
		.DDS1_OutputRelay_s1_write                  (mm_interconnect_0_dds1_outputrelay_s1_write),               //                                     .write
		.DDS1_OutputRelay_s1_readdata               (mm_interconnect_0_dds1_outputrelay_s1_readdata),            //                                     .readdata
		.DDS1_OutputRelay_s1_writedata              (mm_interconnect_0_dds1_outputrelay_s1_writedata),           //                                     .writedata
		.DDS1_OutputRelay_s1_chipselect             (mm_interconnect_0_dds1_outputrelay_s1_chipselect),          //                                     .chipselect
		.DDS1_PhaseOffset_s1_address                (mm_interconnect_0_dds1_phaseoffset_s1_address),             //                  DDS1_PhaseOffset_s1.address
		.DDS1_PhaseOffset_s1_write                  (mm_interconnect_0_dds1_phaseoffset_s1_write),               //                                     .write
		.DDS1_PhaseOffset_s1_readdata               (mm_interconnect_0_dds1_phaseoffset_s1_readdata),            //                                     .readdata
		.DDS1_PhaseOffset_s1_writedata              (mm_interconnect_0_dds1_phaseoffset_s1_writedata),           //                                     .writedata
		.DDS1_PhaseOffset_s1_chipselect             (mm_interconnect_0_dds1_phaseoffset_s1_chipselect),          //                                     .chipselect
		.DDS1_PhaseStep_s1_address                  (mm_interconnect_0_dds1_phasestep_s1_address),               //                    DDS1_PhaseStep_s1.address
		.DDS1_PhaseStep_s1_write                    (mm_interconnect_0_dds1_phasestep_s1_write),                 //                                     .write
		.DDS1_PhaseStep_s1_readdata                 (mm_interconnect_0_dds1_phasestep_s1_readdata),              //                                     .readdata
		.DDS1_PhaseStep_s1_writedata                (mm_interconnect_0_dds1_phasestep_s1_writedata),             //                                     .writedata
		.DDS1_PhaseStep_s1_chipselect               (mm_interconnect_0_dds1_phasestep_s1_chipselect),            //                                     .chipselect
		.DDS1_PM_ModIndex_s1_address                (mm_interconnect_0_dds1_pm_modindex_s1_address),             //                  DDS1_PM_ModIndex_s1.address
		.DDS1_PM_ModIndex_s1_write                  (mm_interconnect_0_dds1_pm_modindex_s1_write),               //                                     .write
		.DDS1_PM_ModIndex_s1_readdata               (mm_interconnect_0_dds1_pm_modindex_s1_readdata),            //                                     .readdata
		.DDS1_PM_ModIndex_s1_writedata              (mm_interconnect_0_dds1_pm_modindex_s1_writedata),           //                                     .writedata
		.DDS1_PM_ModIndex_s1_chipselect             (mm_interconnect_0_dds1_pm_modindex_s1_chipselect),          //                                     .chipselect
		.DDS1_PM_ModPhaseStep_s1_address            (mm_interconnect_0_dds1_pm_modphasestep_s1_address),         //              DDS1_PM_ModPhaseStep_s1.address
		.DDS1_PM_ModPhaseStep_s1_write              (mm_interconnect_0_dds1_pm_modphasestep_s1_write),           //                                     .write
		.DDS1_PM_ModPhaseStep_s1_readdata           (mm_interconnect_0_dds1_pm_modphasestep_s1_readdata),        //                                     .readdata
		.DDS1_PM_ModPhaseStep_s1_writedata          (mm_interconnect_0_dds1_pm_modphasestep_s1_writedata),       //                                     .writedata
		.DDS1_PM_ModPhaseStep_s1_chipselect         (mm_interconnect_0_dds1_pm_modphasestep_s1_chipselect),      //                                     .chipselect
		.DDS1_PWM_Amplitude_s1_address              (mm_interconnect_0_dds1_pwm_amplitude_s1_address),           //                DDS1_PWM_Amplitude_s1.address
		.DDS1_PWM_Amplitude_s1_write                (mm_interconnect_0_dds1_pwm_amplitude_s1_write),             //                                     .write
		.DDS1_PWM_Amplitude_s1_readdata             (mm_interconnect_0_dds1_pwm_amplitude_s1_readdata),          //                                     .readdata
		.DDS1_PWM_Amplitude_s1_writedata            (mm_interconnect_0_dds1_pwm_amplitude_s1_writedata),         //                                     .writedata
		.DDS1_PWM_Amplitude_s1_chipselect           (mm_interconnect_0_dds1_pwm_amplitude_s1_chipselect),        //                                     .chipselect
		.DDS1_PWM_Offset_s1_address                 (mm_interconnect_0_dds1_pwm_offset_s1_address),              //                   DDS1_PWM_Offset_s1.address
		.DDS1_PWM_Offset_s1_write                   (mm_interconnect_0_dds1_pwm_offset_s1_write),                //                                     .write
		.DDS1_PWM_Offset_s1_readdata                (mm_interconnect_0_dds1_pwm_offset_s1_readdata),             //                                     .readdata
		.DDS1_PWM_Offset_s1_writedata               (mm_interconnect_0_dds1_pwm_offset_s1_writedata),            //                                     .writedata
		.DDS1_PWM_Offset_s1_chipselect              (mm_interconnect_0_dds1_pwm_offset_s1_chipselect),           //                                     .chipselect
		.DDS_RESET_s1_address                       (mm_interconnect_0_dds_reset_s1_address),                    //                         DDS_RESET_s1.address
		.DDS_RESET_s1_write                         (mm_interconnect_0_dds_reset_s1_write),                      //                                     .write
		.DDS_RESET_s1_readdata                      (mm_interconnect_0_dds_reset_s1_readdata),                   //                                     .readdata
		.DDS_RESET_s1_writedata                     (mm_interconnect_0_dds_reset_s1_writedata),                  //                                     .writedata
		.DDS_RESET_s1_chipselect                    (mm_interconnect_0_dds_reset_s1_chipselect),                 //                                     .chipselect
		.FLASH_csr_address                          (mm_interconnect_0_flash_csr_address),                       //                            FLASH_csr.address
		.FLASH_csr_write                            (mm_interconnect_0_flash_csr_write),                         //                                     .write
		.FLASH_csr_read                             (mm_interconnect_0_flash_csr_read),                          //                                     .read
		.FLASH_csr_readdata                         (mm_interconnect_0_flash_csr_readdata),                      //                                     .readdata
		.FLASH_csr_writedata                        (mm_interconnect_0_flash_csr_writedata),                     //                                     .writedata
		.FLASH_data_address                         (mm_interconnect_0_flash_data_address),                      //                           FLASH_data.address
		.FLASH_data_write                           (mm_interconnect_0_flash_data_write),                        //                                     .write
		.FLASH_data_read                            (mm_interconnect_0_flash_data_read),                         //                                     .read
		.FLASH_data_readdata                        (mm_interconnect_0_flash_data_readdata),                     //                                     .readdata
		.FLASH_data_writedata                       (mm_interconnect_0_flash_data_writedata),                    //                                     .writedata
		.FLASH_data_burstcount                      (mm_interconnect_0_flash_data_burstcount),                   //                                     .burstcount
		.FLASH_data_readdatavalid                   (mm_interconnect_0_flash_data_readdatavalid),                //                                     .readdatavalid
		.FLASH_data_waitrequest                     (mm_interconnect_0_flash_data_waitrequest),                  //                                     .waitrequest
		.JTAG_UART_avalon_jtag_slave_address        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //          JTAG_UART_avalon_jtag_slave.address
		.JTAG_UART_avalon_jtag_slave_write          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                     .write
		.JTAG_UART_avalon_jtag_slave_read           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                     .read
		.JTAG_UART_avalon_jtag_slave_readdata       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                     .readdata
		.JTAG_UART_avalon_jtag_slave_writedata      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                     .writedata
		.JTAG_UART_avalon_jtag_slave_waitrequest    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                     .waitrequest
		.JTAG_UART_avalon_jtag_slave_chipselect     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                     .chipselect
		.KEYPAD_s1_address                          (mm_interconnect_0_keypad_s1_address),                       //                            KEYPAD_s1.address
		.KEYPAD_s1_write                            (mm_interconnect_0_keypad_s1_write),                         //                                     .write
		.KEYPAD_s1_readdata                         (mm_interconnect_0_keypad_s1_readdata),                      //                                     .readdata
		.KEYPAD_s1_writedata                        (mm_interconnect_0_keypad_s1_writedata),                     //                                     .writedata
		.KEYPAD_s1_chipselect                       (mm_interconnect_0_keypad_s1_chipselect),                    //                                     .chipselect
		.LCD_BackLight_PWM_s1_address               (mm_interconnect_0_lcd_backlight_pwm_s1_address),            //                 LCD_BackLight_PWM_s1.address
		.LCD_BackLight_PWM_s1_write                 (mm_interconnect_0_lcd_backlight_pwm_s1_write),              //                                     .write
		.LCD_BackLight_PWM_s1_readdata              (mm_interconnect_0_lcd_backlight_pwm_s1_readdata),           //                                     .readdata
		.LCD_BackLight_PWM_s1_writedata             (mm_interconnect_0_lcd_backlight_pwm_s1_writedata),          //                                     .writedata
		.LCD_BackLight_PWM_s1_chipselect            (mm_interconnect_0_lcd_backlight_pwm_s1_chipselect),         //                                     .chipselect
		.LCD_Control_s1_address                     (mm_interconnect_0_lcd_control_s1_address),                  //                       LCD_Control_s1.address
		.LCD_Control_s1_write                       (mm_interconnect_0_lcd_control_s1_write),                    //                                     .write
		.LCD_Control_s1_readdata                    (mm_interconnect_0_lcd_control_s1_readdata),                 //                                     .readdata
		.LCD_Control_s1_writedata                   (mm_interconnect_0_lcd_control_s1_writedata),                //                                     .writedata
		.LCD_Control_s1_chipselect                  (mm_interconnect_0_lcd_control_s1_chipselect),               //                                     .chipselect
		.LCD_Data_s1_address                        (mm_interconnect_0_lcd_data_s1_address),                     //                          LCD_Data_s1.address
		.LCD_Data_s1_write                          (mm_interconnect_0_lcd_data_s1_write),                       //                                     .write
		.LCD_Data_s1_readdata                       (mm_interconnect_0_lcd_data_s1_readdata),                    //                                     .readdata
		.LCD_Data_s1_writedata                      (mm_interconnect_0_lcd_data_s1_writedata),                   //                                     .writedata
		.LCD_Data_s1_chipselect                     (mm_interconnect_0_lcd_data_s1_chipselect),                  //                                     .chipselect
		.LCD_DMA_control_port_slave_address         (mm_interconnect_0_lcd_dma_control_port_slave_address),      //           LCD_DMA_control_port_slave.address
		.LCD_DMA_control_port_slave_write           (mm_interconnect_0_lcd_dma_control_port_slave_write),        //                                     .write
		.LCD_DMA_control_port_slave_readdata        (mm_interconnect_0_lcd_dma_control_port_slave_readdata),     //                                     .readdata
		.LCD_DMA_control_port_slave_writedata       (mm_interconnect_0_lcd_dma_control_port_slave_writedata),    //                                     .writedata
		.LCD_DMA_control_port_slave_chipselect      (mm_interconnect_0_lcd_dma_control_port_slave_chipselect),   //                                     .chipselect
		.LOOKUP_RAM_RAM_DDS0_AM_s1_address          (mm_interconnect_0_lookup_ram_ram_dds0_am_s1_address),       //            LOOKUP_RAM_RAM_DDS0_AM_s1.address
		.LOOKUP_RAM_RAM_DDS0_AM_s1_write            (mm_interconnect_0_lookup_ram_ram_dds0_am_s1_write),         //                                     .write
		.LOOKUP_RAM_RAM_DDS0_AM_s1_readdata         (mm_interconnect_0_lookup_ram_ram_dds0_am_s1_readdata),      //                                     .readdata
		.LOOKUP_RAM_RAM_DDS0_AM_s1_writedata        (mm_interconnect_0_lookup_ram_ram_dds0_am_s1_writedata),     //                                     .writedata
		.LOOKUP_RAM_RAM_DDS0_AM_s1_byteenable       (mm_interconnect_0_lookup_ram_ram_dds0_am_s1_byteenable),    //                                     .byteenable
		.LOOKUP_RAM_RAM_DDS0_AM_s1_chipselect       (mm_interconnect_0_lookup_ram_ram_dds0_am_s1_chipselect),    //                                     .chipselect
		.LOOKUP_RAM_RAM_DDS0_AM_s1_clken            (mm_interconnect_0_lookup_ram_ram_dds0_am_s1_clken),         //                                     .clken
		.LOOKUP_RAM_RAM_DDS0_FM_s1_address          (mm_interconnect_0_lookup_ram_ram_dds0_fm_s1_address),       //            LOOKUP_RAM_RAM_DDS0_FM_s1.address
		.LOOKUP_RAM_RAM_DDS0_FM_s1_write            (mm_interconnect_0_lookup_ram_ram_dds0_fm_s1_write),         //                                     .write
		.LOOKUP_RAM_RAM_DDS0_FM_s1_readdata         (mm_interconnect_0_lookup_ram_ram_dds0_fm_s1_readdata),      //                                     .readdata
		.LOOKUP_RAM_RAM_DDS0_FM_s1_writedata        (mm_interconnect_0_lookup_ram_ram_dds0_fm_s1_writedata),     //                                     .writedata
		.LOOKUP_RAM_RAM_DDS0_FM_s1_byteenable       (mm_interconnect_0_lookup_ram_ram_dds0_fm_s1_byteenable),    //                                     .byteenable
		.LOOKUP_RAM_RAM_DDS0_FM_s1_chipselect       (mm_interconnect_0_lookup_ram_ram_dds0_fm_s1_chipselect),    //                                     .chipselect
		.LOOKUP_RAM_RAM_DDS0_FM_s1_clken            (mm_interconnect_0_lookup_ram_ram_dds0_fm_s1_clken),         //                                     .clken
		.LOOKUP_RAM_RAM_DDS0_s1_address             (mm_interconnect_0_lookup_ram_ram_dds0_s1_address),          //               LOOKUP_RAM_RAM_DDS0_s1.address
		.LOOKUP_RAM_RAM_DDS0_s1_write               (mm_interconnect_0_lookup_ram_ram_dds0_s1_write),            //                                     .write
		.LOOKUP_RAM_RAM_DDS0_s1_readdata            (mm_interconnect_0_lookup_ram_ram_dds0_s1_readdata),         //                                     .readdata
		.LOOKUP_RAM_RAM_DDS0_s1_writedata           (mm_interconnect_0_lookup_ram_ram_dds0_s1_writedata),        //                                     .writedata
		.LOOKUP_RAM_RAM_DDS0_s1_byteenable          (mm_interconnect_0_lookup_ram_ram_dds0_s1_byteenable),       //                                     .byteenable
		.LOOKUP_RAM_RAM_DDS0_s1_chipselect          (mm_interconnect_0_lookup_ram_ram_dds0_s1_chipselect),       //                                     .chipselect
		.LOOKUP_RAM_RAM_DDS0_s1_clken               (mm_interconnect_0_lookup_ram_ram_dds0_s1_clken),            //                                     .clken
		.LOOKUP_RAM_RAM_DDS1_AM_s1_address          (mm_interconnect_0_lookup_ram_ram_dds1_am_s1_address),       //            LOOKUP_RAM_RAM_DDS1_AM_s1.address
		.LOOKUP_RAM_RAM_DDS1_AM_s1_write            (mm_interconnect_0_lookup_ram_ram_dds1_am_s1_write),         //                                     .write
		.LOOKUP_RAM_RAM_DDS1_AM_s1_readdata         (mm_interconnect_0_lookup_ram_ram_dds1_am_s1_readdata),      //                                     .readdata
		.LOOKUP_RAM_RAM_DDS1_AM_s1_writedata        (mm_interconnect_0_lookup_ram_ram_dds1_am_s1_writedata),     //                                     .writedata
		.LOOKUP_RAM_RAM_DDS1_AM_s1_byteenable       (mm_interconnect_0_lookup_ram_ram_dds1_am_s1_byteenable),    //                                     .byteenable
		.LOOKUP_RAM_RAM_DDS1_AM_s1_chipselect       (mm_interconnect_0_lookup_ram_ram_dds1_am_s1_chipselect),    //                                     .chipselect
		.LOOKUP_RAM_RAM_DDS1_AM_s1_clken            (mm_interconnect_0_lookup_ram_ram_dds1_am_s1_clken),         //                                     .clken
		.LOOKUP_RAM_RAM_DDS1_FM_s1_address          (mm_interconnect_0_lookup_ram_ram_dds1_fm_s1_address),       //            LOOKUP_RAM_RAM_DDS1_FM_s1.address
		.LOOKUP_RAM_RAM_DDS1_FM_s1_write            (mm_interconnect_0_lookup_ram_ram_dds1_fm_s1_write),         //                                     .write
		.LOOKUP_RAM_RAM_DDS1_FM_s1_readdata         (mm_interconnect_0_lookup_ram_ram_dds1_fm_s1_readdata),      //                                     .readdata
		.LOOKUP_RAM_RAM_DDS1_FM_s1_writedata        (mm_interconnect_0_lookup_ram_ram_dds1_fm_s1_writedata),     //                                     .writedata
		.LOOKUP_RAM_RAM_DDS1_FM_s1_byteenable       (mm_interconnect_0_lookup_ram_ram_dds1_fm_s1_byteenable),    //                                     .byteenable
		.LOOKUP_RAM_RAM_DDS1_FM_s1_chipselect       (mm_interconnect_0_lookup_ram_ram_dds1_fm_s1_chipselect),    //                                     .chipselect
		.LOOKUP_RAM_RAM_DDS1_FM_s1_clken            (mm_interconnect_0_lookup_ram_ram_dds1_fm_s1_clken),         //                                     .clken
		.LOOKUP_RAM_RAM_DDS1_s1_address             (mm_interconnect_0_lookup_ram_ram_dds1_s1_address),          //               LOOKUP_RAM_RAM_DDS1_s1.address
		.LOOKUP_RAM_RAM_DDS1_s1_write               (mm_interconnect_0_lookup_ram_ram_dds1_s1_write),            //                                     .write
		.LOOKUP_RAM_RAM_DDS1_s1_readdata            (mm_interconnect_0_lookup_ram_ram_dds1_s1_readdata),         //                                     .readdata
		.LOOKUP_RAM_RAM_DDS1_s1_writedata           (mm_interconnect_0_lookup_ram_ram_dds1_s1_writedata),        //                                     .writedata
		.LOOKUP_RAM_RAM_DDS1_s1_byteenable          (mm_interconnect_0_lookup_ram_ram_dds1_s1_byteenable),       //                                     .byteenable
		.LOOKUP_RAM_RAM_DDS1_s1_chipselect          (mm_interconnect_0_lookup_ram_ram_dds1_s1_chipselect),       //                                     .chipselect
		.LOOKUP_RAM_RAM_DDS1_s1_clken               (mm_interconnect_0_lookup_ram_ram_dds1_s1_clken),            //                                     .clken
		.LOOKUP_RAM_ISR_s1_address                  (mm_interconnect_0_lookup_ram_isr_s1_address),               //                    LOOKUP_RAM_ISR_s1.address
		.LOOKUP_RAM_ISR_s1_write                    (mm_interconnect_0_lookup_ram_isr_s1_write),                 //                                     .write
		.LOOKUP_RAM_ISR_s1_readdata                 (mm_interconnect_0_lookup_ram_isr_s1_readdata),              //                                     .readdata
		.LOOKUP_RAM_ISR_s1_writedata                (mm_interconnect_0_lookup_ram_isr_s1_writedata),             //                                     .writedata
		.LOOKUP_RAM_ISR_s1_chipselect               (mm_interconnect_0_lookup_ram_isr_s1_chipselect),            //                                     .chipselect
		.NIOS_CPU_debug_mem_slave_address           (mm_interconnect_0_nios_cpu_debug_mem_slave_address),        //             NIOS_CPU_debug_mem_slave.address
		.NIOS_CPU_debug_mem_slave_write             (mm_interconnect_0_nios_cpu_debug_mem_slave_write),          //                                     .write
		.NIOS_CPU_debug_mem_slave_read              (mm_interconnect_0_nios_cpu_debug_mem_slave_read),           //                                     .read
		.NIOS_CPU_debug_mem_slave_readdata          (mm_interconnect_0_nios_cpu_debug_mem_slave_readdata),       //                                     .readdata
		.NIOS_CPU_debug_mem_slave_writedata         (mm_interconnect_0_nios_cpu_debug_mem_slave_writedata),      //                                     .writedata
		.NIOS_CPU_debug_mem_slave_byteenable        (mm_interconnect_0_nios_cpu_debug_mem_slave_byteenable),     //                                     .byteenable
		.NIOS_CPU_debug_mem_slave_waitrequest       (mm_interconnect_0_nios_cpu_debug_mem_slave_waitrequest),    //                                     .waitrequest
		.NIOS_CPU_debug_mem_slave_debugaccess       (mm_interconnect_0_nios_cpu_debug_mem_slave_debugaccess),    //                                     .debugaccess
		.PIO_LED_DEBUG_s1_address                   (mm_interconnect_0_pio_led_debug_s1_address),                //                     PIO_LED_DEBUG_s1.address
		.PIO_LED_DEBUG_s1_write                     (mm_interconnect_0_pio_led_debug_s1_write),                  //                                     .write
		.PIO_LED_DEBUG_s1_readdata                  (mm_interconnect_0_pio_led_debug_s1_readdata),               //                                     .readdata
		.PIO_LED_DEBUG_s1_writedata                 (mm_interconnect_0_pio_led_debug_s1_writedata),              //                                     .writedata
		.PIO_LED_DEBUG_s1_chipselect                (mm_interconnect_0_pio_led_debug_s1_chipselect),             //                                     .chipselect
		.RAM_24K_s1_address                         (mm_interconnect_0_ram_24k_s1_address),                      //                           RAM_24K_s1.address
		.RAM_24K_s1_write                           (mm_interconnect_0_ram_24k_s1_write),                        //                                     .write
		.RAM_24K_s1_readdata                        (mm_interconnect_0_ram_24k_s1_readdata),                     //                                     .readdata
		.RAM_24K_s1_writedata                       (mm_interconnect_0_ram_24k_s1_writedata),                    //                                     .writedata
		.RAM_24K_s1_byteenable                      (mm_interconnect_0_ram_24k_s1_byteenable),                   //                                     .byteenable
		.RAM_24K_s1_chipselect                      (mm_interconnect_0_ram_24k_s1_chipselect),                   //                                     .chipselect
		.RAM_24K_s1_clken                           (mm_interconnect_0_ram_24k_s1_clken),                        //                                     .clken
		.SD_SPI_spi_control_port_address            (mm_interconnect_0_sd_spi_spi_control_port_address),         //              SD_SPI_spi_control_port.address
		.SD_SPI_spi_control_port_write              (mm_interconnect_0_sd_spi_spi_control_port_write),           //                                     .write
		.SD_SPI_spi_control_port_read               (mm_interconnect_0_sd_spi_spi_control_port_read),            //                                     .read
		.SD_SPI_spi_control_port_readdata           (mm_interconnect_0_sd_spi_spi_control_port_readdata),        //                                     .readdata
		.SD_SPI_spi_control_port_writedata          (mm_interconnect_0_sd_spi_spi_control_port_writedata),       //                                     .writedata
		.SD_SPI_spi_control_port_chipselect         (mm_interconnect_0_sd_spi_spi_control_port_chipselect),      //                                     .chipselect
		.SPI_DMA_control_port_slave_address         (mm_interconnect_0_spi_dma_control_port_slave_address),      //           SPI_DMA_control_port_slave.address
		.SPI_DMA_control_port_slave_write           (mm_interconnect_0_spi_dma_control_port_slave_write),        //                                     .write
		.SPI_DMA_control_port_slave_readdata        (mm_interconnect_0_spi_dma_control_port_slave_readdata),     //                                     .readdata
		.SPI_DMA_control_port_slave_writedata       (mm_interconnect_0_spi_dma_control_port_slave_writedata),    //                                     .writedata
		.SPI_DMA_control_port_slave_chipselect      (mm_interconnect_0_spi_dma_control_port_slave_chipselect),   //                                     .chipselect
		.TIMER_DELAY_32bit_s1_address               (mm_interconnect_0_timer_delay_32bit_s1_address),            //                 TIMER_DELAY_32bit_s1.address
		.TIMER_DELAY_32bit_s1_write                 (mm_interconnect_0_timer_delay_32bit_s1_write),              //                                     .write
		.TIMER_DELAY_32bit_s1_readdata              (mm_interconnect_0_timer_delay_32bit_s1_readdata),           //                                     .readdata
		.TIMER_DELAY_32bit_s1_writedata             (mm_interconnect_0_timer_delay_32bit_s1_writedata),          //                                     .writedata
		.TIMER_DELAY_32bit_s1_chipselect            (mm_interconnect_0_timer_delay_32bit_s1_chipselect)          //                                     .chipselect
	);

	NiosII_Processor_irq_mapper irq_mapper (
		.clk           (clk_clk),                  //       clk.clk
		.reset         (cpu_reset),                // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq), // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq), // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq), // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq), // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq), // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq), // receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq), // receiver7.irq
		.receiver8_irq (irq_mapper_receiver8_irq), // receiver8.irq
		.receiver9_irq (irq_mapper_receiver9_irq), // receiver9.irq
		.sender_irq    (nios_cpu_irq_irq)          //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios_cpu_debug_reset_request_reset), // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (cpu_reset),                          // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
