// NiosII_Processor_DDS1.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module NiosII_Processor_DDS1 (
		input  wire        AM_ModIndex_clk_clk,                             //                          AM_ModIndex_clk.clk
		output wire [31:0] AM_ModIndex_external_connection_export,          //          AM_ModIndex_external_connection.export
		input  wire        AM_ModIndex_reset_reset_n,                       //                        AM_ModIndex_reset.reset_n
		input  wire [1:0]  AM_ModIndex_s1_address,                          //                           AM_ModIndex_s1.address
		input  wire        AM_ModIndex_s1_write_n,                          //                                         .write_n
		input  wire [31:0] AM_ModIndex_s1_writedata,                        //                                         .writedata
		input  wire        AM_ModIndex_s1_chipselect,                       //                                         .chipselect
		output wire [31:0] AM_ModIndex_s1_readdata,                         //                                         .readdata
		input  wire        AM_ModPhaseStep_clk_clk,                         //                      AM_ModPhaseStep_clk.clk
		output wire [31:0] AM_ModPhaseStep_external_connection_export,      //      AM_ModPhaseStep_external_connection.export
		input  wire        AM_ModPhaseStep_reset_reset_n,                   //                    AM_ModPhaseStep_reset.reset_n
		input  wire [1:0]  AM_ModPhaseStep_s1_address,                      //                       AM_ModPhaseStep_s1.address
		input  wire        AM_ModPhaseStep_s1_write_n,                      //                                         .write_n
		input  wire [31:0] AM_ModPhaseStep_s1_writedata,                    //                                         .writedata
		input  wire        AM_ModPhaseStep_s1_chipselect,                   //                                         .chipselect
		output wire [31:0] AM_ModPhaseStep_s1_readdata,                     //                                         .readdata
		input  wire        FM_ModDeviationPhase_clk_clk,                    //                 FM_ModDeviationPhase_clk.clk
		output wire [31:0] FM_ModDeviationPhase_external_connection_export, // FM_ModDeviationPhase_external_connection.export
		input  wire        FM_ModDeviationPhase_reset_reset_n,              //               FM_ModDeviationPhase_reset.reset_n
		input  wire [1:0]  FM_ModDeviationPhase_s1_address,                 //                  FM_ModDeviationPhase_s1.address
		input  wire        FM_ModDeviationPhase_s1_write_n,                 //                                         .write_n
		input  wire [31:0] FM_ModDeviationPhase_s1_writedata,               //                                         .writedata
		input  wire        FM_ModDeviationPhase_s1_chipselect,              //                                         .chipselect
		output wire [31:0] FM_ModDeviationPhase_s1_readdata,                //                                         .readdata
		input  wire        FM_ModPhaseStep_clk_clk,                         //                      FM_ModPhaseStep_clk.clk
		output wire [31:0] FM_ModPhaseStep_external_connection_export,      //      FM_ModPhaseStep_external_connection.export
		input  wire        FM_ModPhaseStep_reset_reset_n,                   //                    FM_ModPhaseStep_reset.reset_n
		input  wire [1:0]  FM_ModPhaseStep_s1_address,                      //                       FM_ModPhaseStep_s1.address
		input  wire        FM_ModPhaseStep_s1_write_n,                      //                                         .write_n
		input  wire [31:0] FM_ModPhaseStep_s1_writedata,                    //                                         .writedata
		input  wire        FM_ModPhaseStep_s1_chipselect,                   //                                         .chipselect
		output wire [31:0] FM_ModPhaseStep_s1_readdata,                     //                                         .readdata
		input  wire        OutputRelay_clk_clk,                             //                          OutputRelay_clk.clk
		output wire        OutputRelay_external_connection_export,          //          OutputRelay_external_connection.export
		input  wire        OutputRelay_reset_reset_n,                       //                        OutputRelay_reset.reset_n
		input  wire [1:0]  OutputRelay_s1_address,                          //                           OutputRelay_s1.address
		input  wire        OutputRelay_s1_write_n,                          //                                         .write_n
		input  wire [31:0] OutputRelay_s1_writedata,                        //                                         .writedata
		input  wire        OutputRelay_s1_chipselect,                       //                                         .chipselect
		output wire [31:0] OutputRelay_s1_readdata,                         //                                         .readdata
		input  wire        PM_ModIndex_clk_clk,                             //                          PM_ModIndex_clk.clk
		output wire [31:0] PM_ModIndex_external_connection_export,          //          PM_ModIndex_external_connection.export
		input  wire        PM_ModIndex_reset_reset_n,                       //                        PM_ModIndex_reset.reset_n
		input  wire [1:0]  PM_ModIndex_s1_address,                          //                           PM_ModIndex_s1.address
		input  wire        PM_ModIndex_s1_write_n,                          //                                         .write_n
		input  wire [31:0] PM_ModIndex_s1_writedata,                        //                                         .writedata
		input  wire        PM_ModIndex_s1_chipselect,                       //                                         .chipselect
		output wire [31:0] PM_ModIndex_s1_readdata,                         //                                         .readdata
		input  wire        PM_ModPhaseStep_clk_clk,                         //                      PM_ModPhaseStep_clk.clk
		output wire [31:0] PM_ModPhaseStep_external_connection_export,      //      PM_ModPhaseStep_external_connection.export
		input  wire        PM_ModPhaseStep_reset_reset_n,                   //                    PM_ModPhaseStep_reset.reset_n
		input  wire [1:0]  PM_ModPhaseStep_s1_address,                      //                       PM_ModPhaseStep_s1.address
		input  wire        PM_ModPhaseStep_s1_write_n,                      //                                         .write_n
		input  wire [31:0] PM_ModPhaseStep_s1_writedata,                    //                                         .writedata
		input  wire        PM_ModPhaseStep_s1_chipselect,                   //                                         .chipselect
		output wire [31:0] PM_ModPhaseStep_s1_readdata,                     //                                         .readdata
		input  wire        PWM_Amplitude_clk_clk,                           //                        PWM_Amplitude_clk.clk
		output wire [15:0] PWM_Amplitude_external_connection_export,        //        PWM_Amplitude_external_connection.export
		input  wire        PWM_Amplitude_reset_reset_n,                     //                      PWM_Amplitude_reset.reset_n
		input  wire [1:0]  PWM_Amplitude_s1_address,                        //                         PWM_Amplitude_s1.address
		input  wire        PWM_Amplitude_s1_write_n,                        //                                         .write_n
		input  wire [31:0] PWM_Amplitude_s1_writedata,                      //                                         .writedata
		input  wire        PWM_Amplitude_s1_chipselect,                     //                                         .chipselect
		output wire [31:0] PWM_Amplitude_s1_readdata,                       //                                         .readdata
		input  wire        PWM_Offset_clk_clk,                              //                           PWM_Offset_clk.clk
		output wire [15:0] PWM_Offset_external_connection_export,           //           PWM_Offset_external_connection.export
		input  wire        PWM_Offset_reset_reset_n,                        //                         PWM_Offset_reset.reset_n
		input  wire [1:0]  PWM_Offset_s1_address,                           //                            PWM_Offset_s1.address
		input  wire        PWM_Offset_s1_write_n,                           //                                         .write_n
		input  wire [31:0] PWM_Offset_s1_writedata,                         //                                         .writedata
		input  wire        PWM_Offset_s1_chipselect,                        //                                         .chipselect
		output wire [31:0] PWM_Offset_s1_readdata,                          //                                         .readdata
		input  wire        PhaseOffset_clk_clk,                             //                          PhaseOffset_clk.clk
		output wire [31:0] PhaseOffset_external_connection_export,          //          PhaseOffset_external_connection.export
		input  wire        PhaseOffset_reset_reset_n,                       //                        PhaseOffset_reset.reset_n
		input  wire [1:0]  PhaseOffset_s1_address,                          //                           PhaseOffset_s1.address
		input  wire        PhaseOffset_s1_write_n,                          //                                         .write_n
		input  wire [31:0] PhaseOffset_s1_writedata,                        //                                         .writedata
		input  wire        PhaseOffset_s1_chipselect,                       //                                         .chipselect
		output wire [31:0] PhaseOffset_s1_readdata,                         //                                         .readdata
		input  wire        PhaseStep_clk_clk,                               //                            PhaseStep_clk.clk
		output wire [31:0] PhaseStep_external_connection_export,            //            PhaseStep_external_connection.export
		input  wire        PhaseStep_reset_reset_n,                         //                          PhaseStep_reset.reset_n
		input  wire [1:0]  PhaseStep_s1_address,                            //                             PhaseStep_s1.address
		input  wire        PhaseStep_s1_write_n,                            //                                         .write_n
		input  wire [31:0] PhaseStep_s1_writedata,                          //                                         .writedata
		input  wire        PhaseStep_s1_chipselect,                         //                                         .chipselect
		output wire [31:0] PhaseStep_s1_readdata                            //                                         .readdata
	);

	NiosII_Processor_DDS0_AM_ModIndex am_modindex (
		.clk        (AM_ModIndex_clk_clk),                    //                 clk.clk
		.reset_n    (AM_ModIndex_reset_reset_n),              //               reset.reset_n
		.address    (AM_ModIndex_s1_address),                 //                  s1.address
		.write_n    (AM_ModIndex_s1_write_n),                 //                    .write_n
		.writedata  (AM_ModIndex_s1_writedata),               //                    .writedata
		.chipselect (AM_ModIndex_s1_chipselect),              //                    .chipselect
		.readdata   (AM_ModIndex_s1_readdata),                //                    .readdata
		.out_port   (AM_ModIndex_external_connection_export)  // external_connection.export
	);

	NiosII_Processor_DDS0_AM_ModIndex am_modphasestep (
		.clk        (AM_ModPhaseStep_clk_clk),                    //                 clk.clk
		.reset_n    (AM_ModPhaseStep_reset_reset_n),              //               reset.reset_n
		.address    (AM_ModPhaseStep_s1_address),                 //                  s1.address
		.write_n    (AM_ModPhaseStep_s1_write_n),                 //                    .write_n
		.writedata  (AM_ModPhaseStep_s1_writedata),               //                    .writedata
		.chipselect (AM_ModPhaseStep_s1_chipselect),              //                    .chipselect
		.readdata   (AM_ModPhaseStep_s1_readdata),                //                    .readdata
		.out_port   (AM_ModPhaseStep_external_connection_export)  // external_connection.export
	);

	NiosII_Processor_DDS0_AM_ModIndex fm_moddeviationphase (
		.clk        (FM_ModDeviationPhase_clk_clk),                    //                 clk.clk
		.reset_n    (FM_ModDeviationPhase_reset_reset_n),              //               reset.reset_n
		.address    (FM_ModDeviationPhase_s1_address),                 //                  s1.address
		.write_n    (FM_ModDeviationPhase_s1_write_n),                 //                    .write_n
		.writedata  (FM_ModDeviationPhase_s1_writedata),               //                    .writedata
		.chipselect (FM_ModDeviationPhase_s1_chipselect),              //                    .chipselect
		.readdata   (FM_ModDeviationPhase_s1_readdata),                //                    .readdata
		.out_port   (FM_ModDeviationPhase_external_connection_export)  // external_connection.export
	);

	NiosII_Processor_DDS0_AM_ModIndex fm_modphasestep (
		.clk        (FM_ModPhaseStep_clk_clk),                    //                 clk.clk
		.reset_n    (FM_ModPhaseStep_reset_reset_n),              //               reset.reset_n
		.address    (FM_ModPhaseStep_s1_address),                 //                  s1.address
		.write_n    (FM_ModPhaseStep_s1_write_n),                 //                    .write_n
		.writedata  (FM_ModPhaseStep_s1_writedata),               //                    .writedata
		.chipselect (FM_ModPhaseStep_s1_chipselect),              //                    .chipselect
		.readdata   (FM_ModPhaseStep_s1_readdata),                //                    .readdata
		.out_port   (FM_ModPhaseStep_external_connection_export)  // external_connection.export
	);

	NiosII_Processor_DDS0_OutputRelay outputrelay (
		.clk        (OutputRelay_clk_clk),                    //                 clk.clk
		.reset_n    (OutputRelay_reset_reset_n),              //               reset.reset_n
		.address    (OutputRelay_s1_address),                 //                  s1.address
		.write_n    (OutputRelay_s1_write_n),                 //                    .write_n
		.writedata  (OutputRelay_s1_writedata),               //                    .writedata
		.chipselect (OutputRelay_s1_chipselect),              //                    .chipselect
		.readdata   (OutputRelay_s1_readdata),                //                    .readdata
		.out_port   (OutputRelay_external_connection_export)  // external_connection.export
	);

	NiosII_Processor_DDS0_AM_ModIndex pm_modindex (
		.clk        (PM_ModIndex_clk_clk),                    //                 clk.clk
		.reset_n    (PM_ModIndex_reset_reset_n),              //               reset.reset_n
		.address    (PM_ModIndex_s1_address),                 //                  s1.address
		.write_n    (PM_ModIndex_s1_write_n),                 //                    .write_n
		.writedata  (PM_ModIndex_s1_writedata),               //                    .writedata
		.chipselect (PM_ModIndex_s1_chipselect),              //                    .chipselect
		.readdata   (PM_ModIndex_s1_readdata),                //                    .readdata
		.out_port   (PM_ModIndex_external_connection_export)  // external_connection.export
	);

	NiosII_Processor_DDS0_AM_ModIndex pm_modphasestep (
		.clk        (PM_ModPhaseStep_clk_clk),                    //                 clk.clk
		.reset_n    (PM_ModPhaseStep_reset_reset_n),              //               reset.reset_n
		.address    (PM_ModPhaseStep_s1_address),                 //                  s1.address
		.write_n    (PM_ModPhaseStep_s1_write_n),                 //                    .write_n
		.writedata  (PM_ModPhaseStep_s1_writedata),               //                    .writedata
		.chipselect (PM_ModPhaseStep_s1_chipselect),              //                    .chipselect
		.readdata   (PM_ModPhaseStep_s1_readdata),                //                    .readdata
		.out_port   (PM_ModPhaseStep_external_connection_export)  // external_connection.export
	);

	NiosII_Processor_DDS0_PWM_Amplitude pwm_amplitude (
		.clk        (PWM_Amplitude_clk_clk),                    //                 clk.clk
		.reset_n    (PWM_Amplitude_reset_reset_n),              //               reset.reset_n
		.address    (PWM_Amplitude_s1_address),                 //                  s1.address
		.write_n    (PWM_Amplitude_s1_write_n),                 //                    .write_n
		.writedata  (PWM_Amplitude_s1_writedata),               //                    .writedata
		.chipselect (PWM_Amplitude_s1_chipselect),              //                    .chipselect
		.readdata   (PWM_Amplitude_s1_readdata),                //                    .readdata
		.out_port   (PWM_Amplitude_external_connection_export)  // external_connection.export
	);

	NiosII_Processor_DDS0_PWM_Amplitude pwm_offset (
		.clk        (PWM_Offset_clk_clk),                    //                 clk.clk
		.reset_n    (PWM_Offset_reset_reset_n),              //               reset.reset_n
		.address    (PWM_Offset_s1_address),                 //                  s1.address
		.write_n    (PWM_Offset_s1_write_n),                 //                    .write_n
		.writedata  (PWM_Offset_s1_writedata),               //                    .writedata
		.chipselect (PWM_Offset_s1_chipselect),              //                    .chipselect
		.readdata   (PWM_Offset_s1_readdata),                //                    .readdata
		.out_port   (PWM_Offset_external_connection_export)  // external_connection.export
	);

	NiosII_Processor_DDS0_AM_ModIndex phaseoffset (
		.clk        (PhaseOffset_clk_clk),                    //                 clk.clk
		.reset_n    (PhaseOffset_reset_reset_n),              //               reset.reset_n
		.address    (PhaseOffset_s1_address),                 //                  s1.address
		.write_n    (PhaseOffset_s1_write_n),                 //                    .write_n
		.writedata  (PhaseOffset_s1_writedata),               //                    .writedata
		.chipselect (PhaseOffset_s1_chipselect),              //                    .chipselect
		.readdata   (PhaseOffset_s1_readdata),                //                    .readdata
		.out_port   (PhaseOffset_external_connection_export)  // external_connection.export
	);

	NiosII_Processor_DDS0_AM_ModIndex phasestep (
		.clk        (PhaseStep_clk_clk),                    //                 clk.clk
		.reset_n    (PhaseStep_reset_reset_n),              //               reset.reset_n
		.address    (PhaseStep_s1_address),                 //                  s1.address
		.write_n    (PhaseStep_s1_write_n),                 //                    .write_n
		.writedata  (PhaseStep_s1_writedata),               //                    .writedata
		.chipselect (PhaseStep_s1_chipselect),              //                    .chipselect
		.readdata   (PhaseStep_s1_readdata),                //                    .readdata
		.out_port   (PhaseStep_external_connection_export)  // external_connection.export
	);

endmodule
