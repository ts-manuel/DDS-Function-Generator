// NiosII_Processor_LOOKUP_RAM.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module NiosII_Processor_LOOKUP_RAM (
		input  wire        RAM_DDS0_AM_clk1_clk,            //        RAM_DDS0_AM_clk1.clk
		input  wire        RAM_DDS0_AM_reset1_reset,        //      RAM_DDS0_AM_reset1.reset
		input  wire [9:0]  RAM_DDS0_AM_s1_address,          //          RAM_DDS0_AM_s1.address
		input  wire        RAM_DDS0_AM_s1_clken,            //                        .clken
		input  wire        RAM_DDS0_AM_s1_chipselect,       //                        .chipselect
		input  wire        RAM_DDS0_AM_s1_write,            //                        .write
		output wire [15:0] RAM_DDS0_AM_s1_readdata,         //                        .readdata
		input  wire [15:0] RAM_DDS0_AM_s1_writedata,        //                        .writedata
		input  wire [1:0]  RAM_DDS0_AM_s1_byteenable,       //                        .byteenable
		input  wire [9:0]  RAM_DDS0_AM_s2_address,          //          RAM_DDS0_AM_s2.address
		input  wire        RAM_DDS0_AM_s2_chipselect,       //                        .chipselect
		input  wire        RAM_DDS0_AM_s2_clken,            //                        .clken
		input  wire        RAM_DDS0_AM_s2_write,            //                        .write
		output wire [15:0] RAM_DDS0_AM_s2_readdata,         //                        .readdata
		input  wire [15:0] RAM_DDS0_AM_s2_writedata,        //                        .writedata
		input  wire [1:0]  RAM_DDS0_AM_s2_byteenable,       //                        .byteenable
		input  wire        RAM_DDS0_CLK_in_clk_clk,         //     RAM_DDS0_CLK_in_clk.clk
		input  wire        RAM_DDS0_FM_clk1_clk,            //        RAM_DDS0_FM_clk1.clk
		input  wire        RAM_DDS0_FM_reset1_reset,        //      RAM_DDS0_FM_reset1.reset
		input  wire [9:0]  RAM_DDS0_FM_s1_address,          //          RAM_DDS0_FM_s1.address
		input  wire        RAM_DDS0_FM_s1_clken,            //                        .clken
		input  wire        RAM_DDS0_FM_s1_chipselect,       //                        .chipselect
		input  wire        RAM_DDS0_FM_s1_write,            //                        .write
		output wire [15:0] RAM_DDS0_FM_s1_readdata,         //                        .readdata
		input  wire [15:0] RAM_DDS0_FM_s1_writedata,        //                        .writedata
		input  wire [1:0]  RAM_DDS0_FM_s1_byteenable,       //                        .byteenable
		input  wire [9:0]  RAM_DDS0_FM_s2_address,          //          RAM_DDS0_FM_s2.address
		input  wire        RAM_DDS0_FM_s2_chipselect,       //                        .chipselect
		input  wire        RAM_DDS0_FM_s2_clken,            //                        .clken
		input  wire        RAM_DDS0_FM_s2_write,            //                        .write
		output wire [15:0] RAM_DDS0_FM_s2_readdata,         //                        .readdata
		input  wire [15:0] RAM_DDS0_FM_s2_writedata,        //                        .writedata
		input  wire [1:0]  RAM_DDS0_FM_s2_byteenable,       //                        .byteenable
		input  wire        RAM_DDS0_RESET_in_reset_reset_n, // RAM_DDS0_RESET_in_reset.reset_n
		input  wire        RAM_DDS0_clk1_clk,               //           RAM_DDS0_clk1.clk
		input  wire        RAM_DDS0_reset1_reset,           //         RAM_DDS0_reset1.reset
		input  wire [9:0]  RAM_DDS0_s1_address,             //             RAM_DDS0_s1.address
		input  wire        RAM_DDS0_s1_clken,               //                        .clken
		input  wire        RAM_DDS0_s1_chipselect,          //                        .chipselect
		input  wire        RAM_DDS0_s1_write,               //                        .write
		output wire [15:0] RAM_DDS0_s1_readdata,            //                        .readdata
		input  wire [15:0] RAM_DDS0_s1_writedata,           //                        .writedata
		input  wire [1:0]  RAM_DDS0_s1_byteenable,          //                        .byteenable
		input  wire [9:0]  RAM_DDS0_s2_address,             //             RAM_DDS0_s2.address
		input  wire        RAM_DDS0_s2_chipselect,          //                        .chipselect
		input  wire        RAM_DDS0_s2_clken,               //                        .clken
		input  wire        RAM_DDS0_s2_write,               //                        .write
		output wire [15:0] RAM_DDS0_s2_readdata,            //                        .readdata
		input  wire [15:0] RAM_DDS0_s2_writedata,           //                        .writedata
		input  wire [1:0]  RAM_DDS0_s2_byteenable,          //                        .byteenable
		input  wire        RAM_DDS1_AM_clk1_clk,            //        RAM_DDS1_AM_clk1.clk
		input  wire        RAM_DDS1_AM_reset1_reset,        //      RAM_DDS1_AM_reset1.reset
		input  wire [9:0]  RAM_DDS1_AM_s1_address,          //          RAM_DDS1_AM_s1.address
		input  wire        RAM_DDS1_AM_s1_clken,            //                        .clken
		input  wire        RAM_DDS1_AM_s1_chipselect,       //                        .chipselect
		input  wire        RAM_DDS1_AM_s1_write,            //                        .write
		output wire [15:0] RAM_DDS1_AM_s1_readdata,         //                        .readdata
		input  wire [15:0] RAM_DDS1_AM_s1_writedata,        //                        .writedata
		input  wire [1:0]  RAM_DDS1_AM_s1_byteenable,       //                        .byteenable
		input  wire [9:0]  RAM_DDS1_AM_s2_address,          //          RAM_DDS1_AM_s2.address
		input  wire        RAM_DDS1_AM_s2_chipselect,       //                        .chipselect
		input  wire        RAM_DDS1_AM_s2_clken,            //                        .clken
		input  wire        RAM_DDS1_AM_s2_write,            //                        .write
		output wire [15:0] RAM_DDS1_AM_s2_readdata,         //                        .readdata
		input  wire [15:0] RAM_DDS1_AM_s2_writedata,        //                        .writedata
		input  wire [1:0]  RAM_DDS1_AM_s2_byteenable,       //                        .byteenable
		input  wire        RAM_DDS1_FM_clk1_clk,            //        RAM_DDS1_FM_clk1.clk
		input  wire        RAM_DDS1_FM_reset1_reset,        //      RAM_DDS1_FM_reset1.reset
		input  wire [9:0]  RAM_DDS1_FM_s1_address,          //          RAM_DDS1_FM_s1.address
		input  wire        RAM_DDS1_FM_s1_clken,            //                        .clken
		input  wire        RAM_DDS1_FM_s1_chipselect,       //                        .chipselect
		input  wire        RAM_DDS1_FM_s1_write,            //                        .write
		output wire [15:0] RAM_DDS1_FM_s1_readdata,         //                        .readdata
		input  wire [15:0] RAM_DDS1_FM_s1_writedata,        //                        .writedata
		input  wire [1:0]  RAM_DDS1_FM_s1_byteenable,       //                        .byteenable
		input  wire [9:0]  RAM_DDS1_FM_s2_address,          //          RAM_DDS1_FM_s2.address
		input  wire        RAM_DDS1_FM_s2_chipselect,       //                        .chipselect
		input  wire        RAM_DDS1_FM_s2_clken,            //                        .clken
		input  wire        RAM_DDS1_FM_s2_write,            //                        .write
		output wire [15:0] RAM_DDS1_FM_s2_readdata,         //                        .readdata
		input  wire [15:0] RAM_DDS1_FM_s2_writedata,        //                        .writedata
		input  wire [1:0]  RAM_DDS1_FM_s2_byteenable,       //                        .byteenable
		input  wire        RAM_DDS1_clk1_clk,               //           RAM_DDS1_clk1.clk
		input  wire        RAM_DDS1_reset1_reset,           //         RAM_DDS1_reset1.reset
		input  wire [9:0]  RAM_DDS1_s1_address,             //             RAM_DDS1_s1.address
		input  wire        RAM_DDS1_s1_clken,               //                        .clken
		input  wire        RAM_DDS1_s1_chipselect,          //                        .chipselect
		input  wire        RAM_DDS1_s1_write,               //                        .write
		output wire [15:0] RAM_DDS1_s1_readdata,            //                        .readdata
		input  wire [15:0] RAM_DDS1_s1_writedata,           //                        .writedata
		input  wire [1:0]  RAM_DDS1_s1_byteenable,          //                        .byteenable
		input  wire [9:0]  RAM_DDS1_s2_address,             //             RAM_DDS1_s2.address
		input  wire        RAM_DDS1_s2_chipselect,          //                        .chipselect
		input  wire        RAM_DDS1_s2_clken,               //                        .clken
		input  wire        RAM_DDS1_s2_write,               //                        .write
		output wire [15:0] RAM_DDS1_s2_readdata,            //                        .readdata
		input  wire [15:0] RAM_DDS1_s2_writedata,           //                        .writedata
		input  wire [1:0]  RAM_DDS1_s2_byteenable           //                        .byteenable
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> [RAM_DDS0:reset2, RAM_DDS0_AM:reset2, RAM_DDS0_FM:reset2, RAM_DDS1:reset2, RAM_DDS1_AM:reset2, RAM_DDS1_FM:reset2]

	NiosII_Processor_LOOKUP_RAM_RAM_DDS0 ram_dds0 (
		.clk         (RAM_DDS0_clk1_clk),              //   clk1.clk
		.address     (RAM_DDS0_s1_address),            //     s1.address
		.clken       (RAM_DDS0_s1_clken),              //       .clken
		.chipselect  (RAM_DDS0_s1_chipselect),         //       .chipselect
		.write       (RAM_DDS0_s1_write),              //       .write
		.readdata    (RAM_DDS0_s1_readdata),           //       .readdata
		.writedata   (RAM_DDS0_s1_writedata),          //       .writedata
		.byteenable  (RAM_DDS0_s1_byteenable),         //       .byteenable
		.reset       (RAM_DDS0_reset1_reset),          // reset1.reset
		.address2    (RAM_DDS0_s2_address),            //     s2.address
		.chipselect2 (RAM_DDS0_s2_chipselect),         //       .chipselect
		.clken2      (RAM_DDS0_s2_clken),              //       .clken
		.write2      (RAM_DDS0_s2_write),              //       .write
		.readdata2   (RAM_DDS0_s2_readdata),           //       .readdata
		.writedata2  (RAM_DDS0_s2_writedata),          //       .writedata
		.byteenable2 (RAM_DDS0_s2_byteenable),         //       .byteenable
		.clk2        (RAM_DDS0_CLK_in_clk_clk),        //   clk2.clk
		.reset2      (rst_controller_reset_out_reset), // reset2.reset
		.reset_req   (1'b0),                           // (terminated)
		.freeze      (1'b0),                           // (terminated)
		.reset_req2  (1'b0)                            // (terminated)
	);

	NiosII_Processor_LOOKUP_RAM_RAM_DDS0_AM ram_dds0_am (
		.clk         (RAM_DDS0_AM_clk1_clk),           //   clk1.clk
		.address     (RAM_DDS0_AM_s1_address),         //     s1.address
		.clken       (RAM_DDS0_AM_s1_clken),           //       .clken
		.chipselect  (RAM_DDS0_AM_s1_chipselect),      //       .chipselect
		.write       (RAM_DDS0_AM_s1_write),           //       .write
		.readdata    (RAM_DDS0_AM_s1_readdata),        //       .readdata
		.writedata   (RAM_DDS0_AM_s1_writedata),       //       .writedata
		.byteenable  (RAM_DDS0_AM_s1_byteenable),      //       .byteenable
		.reset       (RAM_DDS0_AM_reset1_reset),       // reset1.reset
		.address2    (RAM_DDS0_AM_s2_address),         //     s2.address
		.chipselect2 (RAM_DDS0_AM_s2_chipselect),      //       .chipselect
		.clken2      (RAM_DDS0_AM_s2_clken),           //       .clken
		.write2      (RAM_DDS0_AM_s2_write),           //       .write
		.readdata2   (RAM_DDS0_AM_s2_readdata),        //       .readdata
		.writedata2  (RAM_DDS0_AM_s2_writedata),       //       .writedata
		.byteenable2 (RAM_DDS0_AM_s2_byteenable),      //       .byteenable
		.clk2        (RAM_DDS0_CLK_in_clk_clk),        //   clk2.clk
		.reset2      (rst_controller_reset_out_reset), // reset2.reset
		.reset_req   (1'b0),                           // (terminated)
		.freeze      (1'b0),                           // (terminated)
		.reset_req2  (1'b0)                            // (terminated)
	);

	NiosII_Processor_LOOKUP_RAM_RAM_DDS0_FM ram_dds0_fm (
		.clk         (RAM_DDS0_FM_clk1_clk),           //   clk1.clk
		.address     (RAM_DDS0_FM_s1_address),         //     s1.address
		.clken       (RAM_DDS0_FM_s1_clken),           //       .clken
		.chipselect  (RAM_DDS0_FM_s1_chipselect),      //       .chipselect
		.write       (RAM_DDS0_FM_s1_write),           //       .write
		.readdata    (RAM_DDS0_FM_s1_readdata),        //       .readdata
		.writedata   (RAM_DDS0_FM_s1_writedata),       //       .writedata
		.byteenable  (RAM_DDS0_FM_s1_byteenable),      //       .byteenable
		.reset       (RAM_DDS0_FM_reset1_reset),       // reset1.reset
		.address2    (RAM_DDS0_FM_s2_address),         //     s2.address
		.chipselect2 (RAM_DDS0_FM_s2_chipselect),      //       .chipselect
		.clken2      (RAM_DDS0_FM_s2_clken),           //       .clken
		.write2      (RAM_DDS0_FM_s2_write),           //       .write
		.readdata2   (RAM_DDS0_FM_s2_readdata),        //       .readdata
		.writedata2  (RAM_DDS0_FM_s2_writedata),       //       .writedata
		.byteenable2 (RAM_DDS0_FM_s2_byteenable),      //       .byteenable
		.clk2        (RAM_DDS0_CLK_in_clk_clk),        //   clk2.clk
		.reset2      (rst_controller_reset_out_reset), // reset2.reset
		.reset_req   (1'b0),                           // (terminated)
		.freeze      (1'b0),                           // (terminated)
		.reset_req2  (1'b0)                            // (terminated)
	);

	NiosII_Processor_LOOKUP_RAM_RAM_DDS1 ram_dds1 (
		.clk         (RAM_DDS1_clk1_clk),              //   clk1.clk
		.address     (RAM_DDS1_s1_address),            //     s1.address
		.clken       (RAM_DDS1_s1_clken),              //       .clken
		.chipselect  (RAM_DDS1_s1_chipselect),         //       .chipselect
		.write       (RAM_DDS1_s1_write),              //       .write
		.readdata    (RAM_DDS1_s1_readdata),           //       .readdata
		.writedata   (RAM_DDS1_s1_writedata),          //       .writedata
		.byteenable  (RAM_DDS1_s1_byteenable),         //       .byteenable
		.reset       (RAM_DDS1_reset1_reset),          // reset1.reset
		.address2    (RAM_DDS1_s2_address),            //     s2.address
		.chipselect2 (RAM_DDS1_s2_chipselect),         //       .chipselect
		.clken2      (RAM_DDS1_s2_clken),              //       .clken
		.write2      (RAM_DDS1_s2_write),              //       .write
		.readdata2   (RAM_DDS1_s2_readdata),           //       .readdata
		.writedata2  (RAM_DDS1_s2_writedata),          //       .writedata
		.byteenable2 (RAM_DDS1_s2_byteenable),         //       .byteenable
		.clk2        (RAM_DDS0_CLK_in_clk_clk),        //   clk2.clk
		.reset2      (rst_controller_reset_out_reset), // reset2.reset
		.reset_req   (1'b0),                           // (terminated)
		.freeze      (1'b0),                           // (terminated)
		.reset_req2  (1'b0)                            // (terminated)
	);

	NiosII_Processor_LOOKUP_RAM_RAM_DDS1_AM ram_dds1_am (
		.clk         (RAM_DDS1_AM_clk1_clk),           //   clk1.clk
		.address     (RAM_DDS1_AM_s1_address),         //     s1.address
		.clken       (RAM_DDS1_AM_s1_clken),           //       .clken
		.chipselect  (RAM_DDS1_AM_s1_chipselect),      //       .chipselect
		.write       (RAM_DDS1_AM_s1_write),           //       .write
		.readdata    (RAM_DDS1_AM_s1_readdata),        //       .readdata
		.writedata   (RAM_DDS1_AM_s1_writedata),       //       .writedata
		.byteenable  (RAM_DDS1_AM_s1_byteenable),      //       .byteenable
		.reset       (RAM_DDS1_AM_reset1_reset),       // reset1.reset
		.address2    (RAM_DDS1_AM_s2_address),         //     s2.address
		.chipselect2 (RAM_DDS1_AM_s2_chipselect),      //       .chipselect
		.clken2      (RAM_DDS1_AM_s2_clken),           //       .clken
		.write2      (RAM_DDS1_AM_s2_write),           //       .write
		.readdata2   (RAM_DDS1_AM_s2_readdata),        //       .readdata
		.writedata2  (RAM_DDS1_AM_s2_writedata),       //       .writedata
		.byteenable2 (RAM_DDS1_AM_s2_byteenable),      //       .byteenable
		.clk2        (RAM_DDS0_CLK_in_clk_clk),        //   clk2.clk
		.reset2      (rst_controller_reset_out_reset), // reset2.reset
		.reset_req   (1'b0),                           // (terminated)
		.freeze      (1'b0),                           // (terminated)
		.reset_req2  (1'b0)                            // (terminated)
	);

	NiosII_Processor_LOOKUP_RAM_RAM_DDS1_FM ram_dds1_fm (
		.clk         (RAM_DDS1_FM_clk1_clk),           //   clk1.clk
		.address     (RAM_DDS1_FM_s1_address),         //     s1.address
		.clken       (RAM_DDS1_FM_s1_clken),           //       .clken
		.chipselect  (RAM_DDS1_FM_s1_chipselect),      //       .chipselect
		.write       (RAM_DDS1_FM_s1_write),           //       .write
		.readdata    (RAM_DDS1_FM_s1_readdata),        //       .readdata
		.writedata   (RAM_DDS1_FM_s1_writedata),       //       .writedata
		.byteenable  (RAM_DDS1_FM_s1_byteenable),      //       .byteenable
		.reset       (RAM_DDS1_FM_reset1_reset),       // reset1.reset
		.address2    (RAM_DDS1_FM_s2_address),         //     s2.address
		.chipselect2 (RAM_DDS1_FM_s2_chipselect),      //       .chipselect
		.clken2      (RAM_DDS1_FM_s2_clken),           //       .clken
		.write2      (RAM_DDS1_FM_s2_write),           //       .write
		.readdata2   (RAM_DDS1_FM_s2_readdata),        //       .readdata
		.writedata2  (RAM_DDS1_FM_s2_writedata),       //       .writedata
		.byteenable2 (RAM_DDS1_FM_s2_byteenable),      //       .byteenable
		.clk2        (RAM_DDS0_CLK_in_clk_clk),        //   clk2.clk
		.reset2      (rst_controller_reset_out_reset), // reset2.reset
		.reset_req   (1'b0),                           // (terminated)
		.freeze      (1'b0),                           // (terminated)
		.reset_req2  (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~RAM_DDS0_RESET_in_reset_reset_n), // reset_in0.reset
		.clk            (RAM_DDS0_CLK_in_clk_clk),          //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),   // reset_out.reset
		.reset_req      (),                                 // (terminated)
		.reset_req_in0  (1'b0),                             // (terminated)
		.reset_in1      (1'b0),                             // (terminated)
		.reset_req_in1  (1'b0),                             // (terminated)
		.reset_in2      (1'b0),                             // (terminated)
		.reset_req_in2  (1'b0),                             // (terminated)
		.reset_in3      (1'b0),                             // (terminated)
		.reset_req_in3  (1'b0),                             // (terminated)
		.reset_in4      (1'b0),                             // (terminated)
		.reset_req_in4  (1'b0),                             // (terminated)
		.reset_in5      (1'b0),                             // (terminated)
		.reset_req_in5  (1'b0),                             // (terminated)
		.reset_in6      (1'b0),                             // (terminated)
		.reset_req_in6  (1'b0),                             // (terminated)
		.reset_in7      (1'b0),                             // (terminated)
		.reset_req_in7  (1'b0),                             // (terminated)
		.reset_in8      (1'b0),                             // (terminated)
		.reset_req_in8  (1'b0),                             // (terminated)
		.reset_in9      (1'b0),                             // (terminated)
		.reset_req_in9  (1'b0),                             // (terminated)
		.reset_in10     (1'b0),                             // (terminated)
		.reset_req_in10 (1'b0),                             // (terminated)
		.reset_in11     (1'b0),                             // (terminated)
		.reset_req_in11 (1'b0),                             // (terminated)
		.reset_in12     (1'b0),                             // (terminated)
		.reset_req_in12 (1'b0),                             // (terminated)
		.reset_in13     (1'b0),                             // (terminated)
		.reset_req_in13 (1'b0),                             // (terminated)
		.reset_in14     (1'b0),                             // (terminated)
		.reset_req_in14 (1'b0),                             // (terminated)
		.reset_in15     (1'b0),                             // (terminated)
		.reset_req_in15 (1'b0)                              // (terminated)
	);

endmodule
